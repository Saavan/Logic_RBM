//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
//
// Create Date: 2019-10-17 17:08:08.996727
// Design Name: vanilla
// Module Name: sigmoidLUT_in6b4p_out16b15p
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 6 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
//
// Additional Comments: Generated by LUT_generator_sigmoid.py
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_in6b4p_out16b15p #(
    parameter PRECISION_INPUT_BITS = 6,
    parameter PRECISION_OUTPUT_BITS = 16
)(
    input[PRECISION_INPUT_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_OUTPUT_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			6'b000000: sigmoid_out <= 16'b0100000000000000;    //sigmoid(0.000000) ≈ 0.500000
			6'b000001: sigmoid_out <= 16'b0100001000000000;    //sigmoid(0.062500) ≈ 0.515625
			6'b000010: sigmoid_out <= 16'b0100001111111111;    //sigmoid(0.125000) ≈ 0.531219
			6'b000011: sigmoid_out <= 16'b0100010111111100;    //sigmoid(0.187500) ≈ 0.546753
			6'b000100: sigmoid_out <= 16'b0100011111110101;    //sigmoid(0.250000) ≈ 0.562164
			6'b000101: sigmoid_out <= 16'b0100100111101011;    //sigmoid(0.312500) ≈ 0.577484
			6'b000110: sigmoid_out <= 16'b0100101111011100;    //sigmoid(0.375000) ≈ 0.592651
			6'b000111: sigmoid_out <= 16'b0100110111001000;    //sigmoid(0.437500) ≈ 0.607666
			6'b001000: sigmoid_out <= 16'b0100111110101101;    //sigmoid(0.500000) ≈ 0.622467
			6'b001001: sigmoid_out <= 16'b0101000110001010;    //sigmoid(0.562500) ≈ 0.637024
			6'b001010: sigmoid_out <= 16'b0101001101100000;    //sigmoid(0.625000) ≈ 0.651367
			6'b001011: sigmoid_out <= 16'b0101010100101100;    //sigmoid(0.687500) ≈ 0.665405
			6'b001100: sigmoid_out <= 16'b0101011011101111;    //sigmoid(0.750000) ≈ 0.679169
			6'b001101: sigmoid_out <= 16'b0101100010101000;    //sigmoid(0.812500) ≈ 0.692627
			6'b001110: sigmoid_out <= 16'b0101101001010111;    //sigmoid(0.875000) ≈ 0.705780
			6'b001111: sigmoid_out <= 16'b0101101111111011;    //sigmoid(0.937500) ≈ 0.718597
			6'b010000: sigmoid_out <= 16'b0101110110010011;    //sigmoid(1.000000) ≈ 0.731049
			6'b010001: sigmoid_out <= 16'b0101111100100000;    //sigmoid(1.062500) ≈ 0.743164
			6'b010010: sigmoid_out <= 16'b0110000010100001;    //sigmoid(1.125000) ≈ 0.754913
			6'b010011: sigmoid_out <= 16'b0110001000010110;    //sigmoid(1.187500) ≈ 0.766296
			6'b010100: sigmoid_out <= 16'b0110001101111111;    //sigmoid(1.250000) ≈ 0.777313
			6'b010101: sigmoid_out <= 16'b0110010011011011;    //sigmoid(1.312500) ≈ 0.787933
			6'b010110: sigmoid_out <= 16'b0110011000101011;    //sigmoid(1.375000) ≈ 0.798187
			6'b010111: sigmoid_out <= 16'b0110011101101111;    //sigmoid(1.437500) ≈ 0.808075
			6'b011000: sigmoid_out <= 16'b0110100010100110;    //sigmoid(1.500000) ≈ 0.817566
			6'b011001: sigmoid_out <= 16'b0110100111010010;    //sigmoid(1.562500) ≈ 0.826721
			6'b011010: sigmoid_out <= 16'b0110101011110001;    //sigmoid(1.625000) ≈ 0.835480
			6'b011011: sigmoid_out <= 16'b0110110000000101;    //sigmoid(1.687500) ≈ 0.843903
			6'b011100: sigmoid_out <= 16'b0110110100001101;    //sigmoid(1.750000) ≈ 0.851959
			6'b011101: sigmoid_out <= 16'b0110111000001001;    //sigmoid(1.812500) ≈ 0.859650
			6'b011110: sigmoid_out <= 16'b0110111011111011;    //sigmoid(1.875000) ≈ 0.867035
			6'b011111: sigmoid_out <= 16'b0110111111100010;    //sigmoid(1.937500) ≈ 0.874084
			6'b100000: sigmoid_out <= 16'b0111000010111110;    //sigmoid(2.000000) ≈ 0.880798
			6'b100001: sigmoid_out <= 16'b0111000110010000;    //sigmoid(2.062500) ≈ 0.887207
			6'b100010: sigmoid_out <= 16'b0111001001011000;    //sigmoid(2.125000) ≈ 0.893311
			6'b100011: sigmoid_out <= 16'b0111001100010110;    //sigmoid(2.187500) ≈ 0.899109
			6'b100100: sigmoid_out <= 16'b0111001111001100;    //sigmoid(2.250000) ≈ 0.904663
			6'b100101: sigmoid_out <= 16'b0111010001111000;    //sigmoid(2.312500) ≈ 0.909912
			6'b100110: sigmoid_out <= 16'b0111010100011011;    //sigmoid(2.375000) ≈ 0.914886
			6'b100111: sigmoid_out <= 16'b0111010110110111;    //sigmoid(2.437500) ≈ 0.919647
			6'b101000: sigmoid_out <= 16'b0111011001001010;    //sigmoid(2.500000) ≈ 0.924133
			6'b101001: sigmoid_out <= 16'b0111011011010110;    //sigmoid(2.562500) ≈ 0.928406
			6'b101010: sigmoid_out <= 16'b0111011101011011;    //sigmoid(2.625000) ≈ 0.932465
			6'b101011: sigmoid_out <= 16'b0111011111011000;    //sigmoid(2.687500) ≈ 0.936279
			6'b101100: sigmoid_out <= 16'b0111100001001111;    //sigmoid(2.750000) ≈ 0.939911
			6'b101101: sigmoid_out <= 16'b0111100011000000;    //sigmoid(2.812500) ≈ 0.943359
			6'b101110: sigmoid_out <= 16'b0111100100101010;    //sigmoid(2.875000) ≈ 0.946594
			6'b101111: sigmoid_out <= 16'b0111100110001111;    //sigmoid(2.937500) ≈ 0.949677
			6'b110000: sigmoid_out <= 16'b0111100111101110;    //sigmoid(3.000000) ≈ 0.952576
			6'b110001: sigmoid_out <= 16'b0111101001001000;    //sigmoid(3.062500) ≈ 0.955322
			6'b110010: sigmoid_out <= 16'b0111101010011101;    //sigmoid(3.125000) ≈ 0.957916
			6'b110011: sigmoid_out <= 16'b0111101011101101;    //sigmoid(3.187500) ≈ 0.960358
			6'b110100: sigmoid_out <= 16'b0111101100111001;    //sigmoid(3.250000) ≈ 0.962677
			6'b110101: sigmoid_out <= 16'b0111101110000000;    //sigmoid(3.312500) ≈ 0.964844
			6'b110110: sigmoid_out <= 16'b0111101111000100;    //sigmoid(3.375000) ≈ 0.966919
			6'b110111: sigmoid_out <= 16'b0111110000000011;    //sigmoid(3.437500) ≈ 0.968842
			6'b111000: sigmoid_out <= 16'b0111110000111111;    //sigmoid(3.500000) ≈ 0.970673
			6'b111001: sigmoid_out <= 16'b0111110001111000;    //sigmoid(3.562500) ≈ 0.972412
			6'b111010: sigmoid_out <= 16'b0111110010101101;    //sigmoid(3.625000) ≈ 0.974030
			6'b111011: sigmoid_out <= 16'b0111110011100000;    //sigmoid(3.687500) ≈ 0.975586
			6'b111100: sigmoid_out <= 16'b0111110100001111;    //sigmoid(3.750000) ≈ 0.977020
			6'b111101: sigmoid_out <= 16'b0111110100111100;    //sigmoid(3.812500) ≈ 0.978394
			6'b111110: sigmoid_out <= 16'b0111110101100110;    //sigmoid(3.875000) ≈ 0.979675
			6'b111111: sigmoid_out <= 16'b0111110110001101;    //sigmoid(3.937500) ≈ 0.980865

        endcase
    end
endmodule