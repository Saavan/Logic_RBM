//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
//
// Create Date: 2019-07-05 14:50:01.745601
// Design Name: vanilla
// Module Name: sigmoidLUT_in8b4p_out32b31p
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 8 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
//
// Additional Comments: Generated by LUT_generator_sigmoid.py
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_in8b4p_out32b31p #(
    parameter PRECISION_INPUT_BITS = 8,
    parameter PRECISION_OUTPUT_BITS = 32
)(
    input[PRECISION_INPUT_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_OUTPUT_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			8'b00000000: sigmoid_out <= 32'b01000000000000000000000000000000;    //sigmoid(0.000000) ≈ 0.500000
			8'b00000001: sigmoid_out <= 32'b01000001111111111101010101011010;    //sigmoid(0.062500) ≈ 0.515620
			8'b00000010: sigmoid_out <= 32'b01000011111111101010101100110011;    //sigmoid(0.125000) ≈ 0.531209
			8'b00000011: sigmoid_out <= 32'b01000101111110111000010000001001;    //sigmoid(0.187500) ≈ 0.546738
			8'b00000100: sigmoid_out <= 32'b01000111111101010110011001001011;    //sigmoid(0.250000) ≈ 0.562177
			8'b00000101: sigmoid_out <= 32'b01001001111010110101111000111110;    //sigmoid(0.312500) ≈ 0.577495
			8'b00000110: sigmoid_out <= 32'b01001011110111000111111111001000;    //sigmoid(0.375000) ≈ 0.592667
			8'b00000111: sigmoid_out <= 32'b01001101110001111110100000100001;    //sigmoid(0.437500) ≈ 0.607663
			8'b00001000: sigmoid_out <= 32'b01001111101011001011111101010011;    //sigmoid(0.500000) ≈ 0.622459
			8'b00001001: sigmoid_out <= 32'b01010001100010100011100110011110;    //sigmoid(0.562500) ≈ 0.637031
			8'b00001010: sigmoid_out <= 32'b01010011010111111001100010100001;    //sigmoid(0.625000) ≈ 0.651355
			8'b00001011: sigmoid_out <= 32'b01010101001011000010110001010110;    //sigmoid(0.687500) ≈ 0.665411
			8'b00001100: sigmoid_out <= 32'b01010110111011110101001111011111;    //sigmoid(0.750000) ≈ 0.679179
			8'b00001101: sigmoid_out <= 32'b01011000101010000111111000010101;    //sigmoid(0.812500) ≈ 0.692642
			8'b00001110: sigmoid_out <= 32'b01011010010101110010100111101110;    //sigmoid(0.875000) ≈ 0.705785
			8'b00001111: sigmoid_out <= 32'b01011011111110101110011010101100;    //sigmoid(0.937500) ≈ 0.718594
			8'b00010000: sigmoid_out <= 32'b01011101100100110101001111010111;    //sigmoid(1.000000) ≈ 0.731059
			8'b00010001: sigmoid_out <= 32'b01011111001000000010000100011010;    //sigmoid(1.062500) ≈ 0.743168
			8'b00010010: sigmoid_out <= 32'b01100000101000010000110111100110;    //sigmoid(1.125000) ≈ 0.754915
			8'b00010011: sigmoid_out <= 32'b01100010000101011110100011111100;    //sigmoid(1.187500) ≈ 0.766294
			8'b00010100: sigmoid_out <= 32'b01100011011111101000111111010101;    //sigmoid(1.250000) ≈ 0.777300
			8'b00010101: sigmoid_out <= 32'b01100100110110101110110111101110;    //sigmoid(1.312500) ≈ 0.787931
			8'b00010110: sigmoid_out <= 32'b01100110001010101111101111111101;    //sigmoid(1.375000) ≈ 0.798187
			8'b00010111: sigmoid_out <= 32'b01100111011011101011111100011000;    //sigmoid(1.437500) ≈ 0.808067
			8'b00011000: sigmoid_out <= 32'b01101000101001100100011111001011;    //sigmoid(1.500000) ≈ 0.817574
			8'b00011001: sigmoid_out <= 32'b01101001110100011011000100101011;    //sigmoid(1.562500) ≈ 0.826712
			8'b00011010: sigmoid_out <= 32'b01101010111100010001111111100010;    //sigmoid(1.625000) ≈ 0.835484
			8'b00011011: sigmoid_out <= 32'b01101100000001001100000100110101;    //sigmoid(1.687500) ≈ 0.843895
			8'b00011100: sigmoid_out <= 32'b01101101000011001100101000010111;    //sigmoid(1.750000) ≈ 0.851953
			8'b00011101: sigmoid_out <= 32'b01101110000010010111011000110111;    //sigmoid(1.812500) ≈ 0.859664
			8'b00011110: sigmoid_out <= 32'b01101110111110110000011100011100;    //sigmoid(1.875000) ≈ 0.867036
			8'b00011111: sigmoid_out <= 32'b01101111111000011100001101001010;    //sigmoid(1.937500) ≈ 0.874077
			8'b00100000: sigmoid_out <= 32'b01110000101111011111010101101010;    //sigmoid(2.000000) ≈ 0.880797
			8'b00100001: sigmoid_out <= 32'b01110001100011111110101110001101;    //sigmoid(2.062500) ≈ 0.887205
			8'b00100010: sigmoid_out <= 32'b01110010010101111111011001101110;    //sigmoid(2.125000) ≈ 0.893309
			8'b00100011: sigmoid_out <= 32'b01110011000101100110100011000111;    //sigmoid(2.187500) ≈ 0.899121
			8'b00100100: sigmoid_out <= 32'b01110011110010111001011010110111;    //sigmoid(2.250000) ≈ 0.904651
			8'b00100101: sigmoid_out <= 32'b01110100011101111101010100110001;    //sigmoid(2.312500) ≈ 0.909907
			8'b00100110: sigmoid_out <= 32'b01110101000110110111100101111000;    //sigmoid(2.375000) ≈ 0.914901
			8'b00100111: sigmoid_out <= 32'b01110101101101101101100010110010;    //sigmoid(2.437500) ≈ 0.919643
			8'b00101000: sigmoid_out <= 32'b01110110010010100100011101110111;    //sigmoid(2.500000) ≈ 0.924142
			8'b00101001: sigmoid_out <= 32'b01110110110101100001100101111110;    //sigmoid(2.562500) ≈ 0.928409
			8'b00101010: sigmoid_out <= 32'b01110111010110101010000101001001;    //sigmoid(2.625000) ≈ 0.932453
			8'b00101011: sigmoid_out <= 32'b01110111110110000010111111100100;    //sigmoid(2.687500) ≈ 0.936285
			8'b00101100: sigmoid_out <= 32'b01111000010011110001010010100101;    //sigmoid(2.750000) ≈ 0.939913
			8'b00101101: sigmoid_out <= 32'b01111000101111111001110100000011;    //sigmoid(2.812500) ≈ 0.943348
			8'b00101110: sigmoid_out <= 32'b01111001001010100001010001100111;    //sigmoid(2.875000) ≈ 0.946597
			8'b00101111: sigmoid_out <= 32'b01111001100011101100010000001110;    //sigmoid(2.937500) ≈ 0.949669
			8'b00110000: sigmoid_out <= 32'b01111001111011011111001011110001;    //sigmoid(3.000000) ≈ 0.952574
			8'b00110001: sigmoid_out <= 32'b01111010010001111110010110110010;    //sigmoid(3.062500) ≈ 0.955319
			8'b00110010: sigmoid_out <= 32'b01111010100111001101111010001101;    //sigmoid(3.125000) ≈ 0.957912
			8'b00110011: sigmoid_out <= 32'b01111010111011010001110101010001;    //sigmoid(3.187500) ≈ 0.960361
			8'b00110100: sigmoid_out <= 32'b01111011001110001101111101100000;    //sigmoid(3.250000) ≈ 0.962673
			8'b00110101: sigmoid_out <= 32'b01111011100000000101111110101001;    //sigmoid(3.312500) ≈ 0.964855
			8'b00110110: sigmoid_out <= 32'b01111011110000111101011010110010;    //sigmoid(3.375000) ≈ 0.966914
			8'b00110111: sigmoid_out <= 32'b01111100000000110111101010011101;    //sigmoid(3.437500) ≈ 0.968856
			8'b00111000: sigmoid_out <= 32'b01111100001111110111111100110000;    //sigmoid(3.500000) ≈ 0.970688
			8'b00111001: sigmoid_out <= 32'b01111100011110000001010111100001;    //sigmoid(3.562500) ≈ 0.972415
			8'b00111010: sigmoid_out <= 32'b01111100101011010110110111101000;    //sigmoid(3.625000) ≈ 0.974043
			8'b00111011: sigmoid_out <= 32'b01111100110111111011010001000101;    //sigmoid(3.687500) ≈ 0.975577
			8'b00111100: sigmoid_out <= 32'b01111101000011110001001111011010;    //sigmoid(3.750000) ≈ 0.977023
			8'b00111101: sigmoid_out <= 32'b01111101001110111011010101110010;    //sigmoid(3.812500) ≈ 0.978385
			8'b00111110: sigmoid_out <= 32'b01111101011001011011111111011100;    //sigmoid(3.875000) ≈ 0.979668
			8'b00111111: sigmoid_out <= 32'b01111101100011010101011111110100;    //sigmoid(3.937500) ≈ 0.980876
			8'b01000000: sigmoid_out <= 32'b01111101101100101010000010111100;    //sigmoid(4.000000) ≈ 0.982014
			8'b01000001: sigmoid_out <= 32'b01111101110101011011101101101100;    //sigmoid(4.062500) ≈ 0.983085
			8'b01000010: sigmoid_out <= 32'b01111101111101101100011110000100;    //sigmoid(4.125000) ≈ 0.984094
			8'b01000011: sigmoid_out <= 32'b01111110000101011110001011011101;    //sigmoid(4.187500) ≈ 0.985043
			8'b01000100: sigmoid_out <= 32'b01111110001100110010100110111111;    //sigmoid(4.250000) ≈ 0.985936
			8'b01000101: sigmoid_out <= 32'b01111110010011101011011011101111;    //sigmoid(4.312500) ≈ 0.986777
			8'b01000110: sigmoid_out <= 32'b01111110011010001010001111000001;    //sigmoid(4.375000) ≈ 0.987568
			8'b01000111: sigmoid_out <= 32'b01111110100000010000100000101101;    //sigmoid(4.437500) ≈ 0.988313
			8'b01001000: sigmoid_out <= 32'b01111110100101111111101011011000;    //sigmoid(4.500000) ≈ 0.989013
			8'b01001001: sigmoid_out <= 32'b01111110101011011001000100101101;    //sigmoid(4.562500) ≈ 0.989672
			8'b01001010: sigmoid_out <= 32'b01111110110000011101111101100110;    //sigmoid(4.625000) ≈ 0.990292
			8'b01001011: sigmoid_out <= 32'b01111110110101001111100010011011;    //sigmoid(4.687500) ≈ 0.990874
			8'b01001100: sigmoid_out <= 32'b01111110111001101110111011010110;    //sigmoid(4.750000) ≈ 0.991423
			8'b01001101: sigmoid_out <= 32'b01111110111101111101001100011101;    //sigmoid(4.812500) ≈ 0.991938
			8'b01001110: sigmoid_out <= 32'b01111111000001111011010101111110;    //sigmoid(4.875000) ≈ 0.992423
			8'b01001111: sigmoid_out <= 32'b01111111000101101010010100100000;    //sigmoid(4.937500) ≈ 0.992879
			8'b01010000: sigmoid_out <= 32'b01111111001001001011000001001100;    //sigmoid(5.000000) ≈ 0.993307
			8'b01010001: sigmoid_out <= 32'b01111111001100011110010001111010;    //sigmoid(5.062500) ≈ 0.993710
			8'b01010010: sigmoid_out <= 32'b01111111001111100100111001011100;    //sigmoid(5.125000) ≈ 0.994089
			8'b01010011: sigmoid_out <= 32'b01111111010010011111100111101010;    //sigmoid(5.187500) ≈ 0.994445
			8'b01010100: sigmoid_out <= 32'b01111111010101001111001001101001;    //sigmoid(5.250000) ≈ 0.994780
			8'b01010101: sigmoid_out <= 32'b01111111010111110100001001111001;    //sigmoid(5.312500) ≈ 0.995095
			8'b01010110: sigmoid_out <= 32'b01111111011010001111010000011011;    //sigmoid(5.375000) ≈ 0.995390
			8'b01010111: sigmoid_out <= 32'b01111111011100100001000010111010;    //sigmoid(5.437500) ≈ 0.995668
			8'b01011000: sigmoid_out <= 32'b01111111011110101010000100110110;    //sigmoid(5.500000) ≈ 0.995930
			8'b01011001: sigmoid_out <= 32'b01111111100000101010110111101000;    //sigmoid(5.562500) ≈ 0.996176
			8'b01011010: sigmoid_out <= 32'b01111111100010100011111010101101;    //sigmoid(5.625000) ≈ 0.996406
			8'b01011011: sigmoid_out <= 32'b01111111100100010101101011101100;    //sigmoid(5.687500) ≈ 0.996623
			8'b01011100: sigmoid_out <= 32'b01111111100110000000100110011011;    //sigmoid(5.750000) ≈ 0.996827
			8'b01011101: sigmoid_out <= 32'b01111111100111100101000101001001;    //sigmoid(5.812500) ≈ 0.997019
			8'b01011110: sigmoid_out <= 32'b01111111101001000011100000011111;    //sigmoid(5.875000) ≈ 0.997199
			8'b01011111: sigmoid_out <= 32'b01111111101010011100001111101011;    //sigmoid(5.937500) ≈ 0.997368
			8'b01100000: sigmoid_out <= 32'b01111111101011101111101000100010;    //sigmoid(6.000000) ≈ 0.997527
			8'b01100001: sigmoid_out <= 32'b01111111101100111101111111100110;    //sigmoid(6.062500) ≈ 0.997677
			8'b01100010: sigmoid_out <= 32'b01111111101110000111101000001100;    //sigmoid(6.125000) ≈ 0.997817
			8'b01100011: sigmoid_out <= 32'b01111111101111001100110100011110;    //sigmoid(6.187500) ≈ 0.997949
			8'b01100100: sigmoid_out <= 32'b01111111110000001101110101100001;    //sigmoid(6.250000) ≈ 0.998073
			8'b01100101: sigmoid_out <= 32'b01111111110001001010111011011001;    //sigmoid(6.312500) ≈ 0.998190
			8'b01100110: sigmoid_out <= 32'b01111111110010000100010101001110;    //sigmoid(6.375000) ≈ 0.998299
			8'b01100111: sigmoid_out <= 32'b01111111110010111010010001001101;    //sigmoid(6.437500) ≈ 0.998402
			8'b01101000: sigmoid_out <= 32'b01111111110011101100111100101100;    //sigmoid(6.500000) ≈ 0.998499
			8'b01101001: sigmoid_out <= 32'b01111111110100011100100100001110;    //sigmoid(6.562500) ≈ 0.998590
			8'b01101010: sigmoid_out <= 32'b01111111110101001001010011101000;    //sigmoid(6.625000) ≈ 0.998675
			8'b01101011: sigmoid_out <= 32'b01111111110101110011010101111111;    //sigmoid(6.687500) ≈ 0.998755
			8'b01101100: sigmoid_out <= 32'b01111111110110011010110101110000;    //sigmoid(6.750000) ≈ 0.998830
			8'b01101101: sigmoid_out <= 32'b01111111110110111111111100101101;    //sigmoid(6.812500) ≈ 0.998901
			8'b01101110: sigmoid_out <= 32'b01111111110111100010110100000101;    //sigmoid(6.875000) ≈ 0.998968
			8'b01101111: sigmoid_out <= 32'b01111111111000000011100100100010;    //sigmoid(6.937500) ≈ 0.999030
			8'b01110000: sigmoid_out <= 32'b01111111111000100010010110001100;    //sigmoid(7.000000) ≈ 0.999089
			8'b01110001: sigmoid_out <= 32'b01111111111000111111010000101111;    //sigmoid(7.062500) ≈ 0.999144
			8'b01110010: sigmoid_out <= 32'b01111111111001011010011011010111;    //sigmoid(7.125000) ≈ 0.999196
			8'b01110011: sigmoid_out <= 32'b01111111111001110011111100110011;    //sigmoid(7.187500) ≈ 0.999245
			8'b01110100: sigmoid_out <= 32'b01111111111010001011111011011010;    //sigmoid(7.250000) ≈ 0.999290
			8'b01110101: sigmoid_out <= 32'b01111111111010100010011101001100;    //sigmoid(7.312500) ≈ 0.999333
			8'b01110110: sigmoid_out <= 32'b01111111111010110111100111101110;    //sigmoid(7.375000) ≈ 0.999374
			8'b01110111: sigmoid_out <= 32'b01111111111011001011100000010010;    //sigmoid(7.437500) ≈ 0.999412
			8'b01111000: sigmoid_out <= 32'b01111111111011011110001011110101;    //sigmoid(7.500000) ≈ 0.999447
			8'b01111001: sigmoid_out <= 32'b01111111111011101111101111000001;    //sigmoid(7.562500) ≈ 0.999481
			8'b01111010: sigmoid_out <= 32'b01111111111100000000001110001111;    //sigmoid(7.625000) ≈ 0.999512
			8'b01111011: sigmoid_out <= 32'b01111111111100001111101101100101;    //sigmoid(7.687500) ≈ 0.999542
			8'b01111100: sigmoid_out <= 32'b01111111111100011110010000111010;    //sigmoid(7.750000) ≈ 0.999569
			8'b01111101: sigmoid_out <= 32'b01111111111100101011111011110111;    //sigmoid(7.812500) ≈ 0.999596
			8'b01111110: sigmoid_out <= 32'b01111111111100111000110001110101;    //sigmoid(7.875000) ≈ 0.999620
			8'b01111111: sigmoid_out <= 32'b01111111111101000100110110000011;    //sigmoid(7.937500) ≈ 0.999643
			8'b10000000: sigmoid_out <= 32'b01111111111101010000001011100001;    //sigmoid(8.000000) ≈ 0.999665
			8'b10000001: sigmoid_out <= 32'b01111111111101011010110101000100;    //sigmoid(8.062500) ≈ 0.999685
			8'b10000010: sigmoid_out <= 32'b01111111111101100100110101010101;    //sigmoid(8.125000) ≈ 0.999704
			8'b10000011: sigmoid_out <= 32'b01111111111101101110001110110101;    //sigmoid(8.187500) ≈ 0.999722
			8'b10000100: sigmoid_out <= 32'b01111111111101110111000011111010;    //sigmoid(8.250000) ≈ 0.999739
			8'b10000101: sigmoid_out <= 32'b01111111111101111111010110110001;    //sigmoid(8.312500) ≈ 0.999755
			8'b10000110: sigmoid_out <= 32'b01111111111110000111001001011111;    //sigmoid(8.375000) ≈ 0.999769
			8'b10000111: sigmoid_out <= 32'b01111111111110001110011101111111;    //sigmoid(8.437500) ≈ 0.999783
			8'b10001000: sigmoid_out <= 32'b01111111111110010101010110001000;    //sigmoid(8.500000) ≈ 0.999797
			8'b10001001: sigmoid_out <= 32'b01111111111110011011110011100111;    //sigmoid(8.562500) ≈ 0.999809
			8'b10001010: sigmoid_out <= 32'b01111111111110100001111000000011;    //sigmoid(8.625000) ≈ 0.999820
			8'b10001011: sigmoid_out <= 32'b01111111111110100111100100111101;    //sigmoid(8.687500) ≈ 0.999831
			8'b10001100: sigmoid_out <= 32'b01111111111110101100111011110001;    //sigmoid(8.750000) ≈ 0.999842
			8'b10001101: sigmoid_out <= 32'b01111111111110110001111101110100;    //sigmoid(8.812500) ≈ 0.999851
			8'b10001110: sigmoid_out <= 32'b01111111111110110110101100010110;    //sigmoid(8.875000) ≈ 0.999860
			8'b10001111: sigmoid_out <= 32'b01111111111110111011001000100100;    //sigmoid(8.937500) ≈ 0.999869
			8'b10010000: sigmoid_out <= 32'b01111111111110111111010011100100;    //sigmoid(9.000000) ≈ 0.999877
			8'b10010001: sigmoid_out <= 32'b01111111111111000011001110011001;    //sigmoid(9.062500) ≈ 0.999884
			8'b10010010: sigmoid_out <= 32'b01111111111111000110111010000010;    //sigmoid(9.125000) ≈ 0.999891
			8'b10010011: sigmoid_out <= 32'b01111111111111001010010111011001;    //sigmoid(9.187500) ≈ 0.999898
			8'b10010100: sigmoid_out <= 32'b01111111111111001101100111010110;    //sigmoid(9.250000) ≈ 0.999904
			8'b10010101: sigmoid_out <= 32'b01111111111111010000101010101100;    //sigmoid(9.312500) ≈ 0.999910
			8'b10010110: sigmoid_out <= 32'b01111111111111010011100010001110;    //sigmoid(9.375000) ≈ 0.999915
			8'b10010111: sigmoid_out <= 32'b01111111111111010110001110101000;    //sigmoid(9.437500) ≈ 0.999920
			8'b10011000: sigmoid_out <= 32'b01111111111111011000110000100101;    //sigmoid(9.500000) ≈ 0.999925
			8'b10011001: sigmoid_out <= 32'b01111111111111011011001000101110;    //sigmoid(9.562500) ≈ 0.999930
			8'b10011010: sigmoid_out <= 32'b01111111111111011101010111101010;    //sigmoid(9.625000) ≈ 0.999934
			8'b10011011: sigmoid_out <= 32'b01111111111111011111011101111100;    //sigmoid(9.687500) ≈ 0.999938
			8'b10011100: sigmoid_out <= 32'b01111111111111100001011100000100;    //sigmoid(9.750000) ≈ 0.999942
			8'b10011101: sigmoid_out <= 32'b01111111111111100011010010100100;    //sigmoid(9.812500) ≈ 0.999945
			8'b10011110: sigmoid_out <= 32'b01111111111111100101000001111001;    //sigmoid(9.875000) ≈ 0.999949
			8'b10011111: sigmoid_out <= 32'b01111111111111100110101010011101;    //sigmoid(9.937500) ≈ 0.999952
			8'b10100000: sigmoid_out <= 32'b01111111111111101000001100101101;    //sigmoid(10.000000) ≈ 0.999955
			8'b10100001: sigmoid_out <= 32'b01111111111111101001101000111111;    //sigmoid(10.062500) ≈ 0.999957
			8'b10100010: sigmoid_out <= 32'b01111111111111101010111111101100;    //sigmoid(10.125000) ≈ 0.999960
			8'b10100011: sigmoid_out <= 32'b01111111111111101100010001001000;    //sigmoid(10.187500) ≈ 0.999962
			8'b10100100: sigmoid_out <= 32'b01111111111111101101011101101001;    //sigmoid(10.250000) ≈ 0.999965
			8'b10100101: sigmoid_out <= 32'b01111111111111101110100101100001;    //sigmoid(10.312500) ≈ 0.999967
			8'b10100110: sigmoid_out <= 32'b01111111111111101111101001000010;    //sigmoid(10.375000) ≈ 0.999969
			8'b10100111: sigmoid_out <= 32'b01111111111111110000101000011110;    //sigmoid(10.437500) ≈ 0.999971
			8'b10101000: sigmoid_out <= 32'b01111111111111110001100100000100;    //sigmoid(10.500000) ≈ 0.999972
			8'b10101001: sigmoid_out <= 32'b01111111111111110010011100000010;    //sigmoid(10.562500) ≈ 0.999974
			8'b10101010: sigmoid_out <= 32'b01111111111111110011010000101000;    //sigmoid(10.625000) ≈ 0.999976
			8'b10101011: sigmoid_out <= 32'b01111111111111110100000010000001;    //sigmoid(10.687500) ≈ 0.999977
			8'b10101100: sigmoid_out <= 32'b01111111111111110100110000011011;    //sigmoid(10.750000) ≈ 0.999979
			8'b10101101: sigmoid_out <= 32'b01111111111111110101011100000001;    //sigmoid(10.812500) ≈ 0.999980
			8'b10101110: sigmoid_out <= 32'b01111111111111110110000100111111;    //sigmoid(10.875000) ≈ 0.999981
			8'b10101111: sigmoid_out <= 32'b01111111111111110110101011011101;    //sigmoid(10.937500) ≈ 0.999982
			8'b10110000: sigmoid_out <= 32'b01111111111111110111001111100110;    //sigmoid(11.000000) ≈ 0.999983
			8'b10110001: sigmoid_out <= 32'b01111111111111110111110001100011;    //sigmoid(11.062500) ≈ 0.999984
			8'b10110010: sigmoid_out <= 32'b01111111111111111000010001011100;    //sigmoid(11.125000) ≈ 0.999985
			8'b10110011: sigmoid_out <= 32'b01111111111111111000101111011010;    //sigmoid(11.187500) ≈ 0.999986
			8'b10110100: sigmoid_out <= 32'b01111111111111111001001011100011;    //sigmoid(11.250000) ≈ 0.999987
			8'b10110101: sigmoid_out <= 32'b01111111111111111001100110000000;    //sigmoid(11.312500) ≈ 0.999988
			8'b10110110: sigmoid_out <= 32'b01111111111111111001111110110110;    //sigmoid(11.375000) ≈ 0.999989
			8'b10110111: sigmoid_out <= 32'b01111111111111111010010110001011;    //sigmoid(11.437500) ≈ 0.999989
			8'b10111000: sigmoid_out <= 32'b01111111111111111010101100000110;    //sigmoid(11.500000) ≈ 0.999990
			8'b10111001: sigmoid_out <= 32'b01111111111111111011000000101100;    //sigmoid(11.562500) ≈ 0.999990
			8'b10111010: sigmoid_out <= 32'b01111111111111111011010100000010;    //sigmoid(11.625000) ≈ 0.999991
			8'b10111011: sigmoid_out <= 32'b01111111111111111011100110001101;    //sigmoid(11.687500) ≈ 0.999992
			8'b10111100: sigmoid_out <= 32'b01111111111111111011110111010010;    //sigmoid(11.750000) ≈ 0.999992
			8'b10111101: sigmoid_out <= 32'b01111111111111111100000111010100;    //sigmoid(11.812500) ≈ 0.999993
			8'b10111110: sigmoid_out <= 32'b01111111111111111100010110011001;    //sigmoid(11.875000) ≈ 0.999993
			8'b10111111: sigmoid_out <= 32'b01111111111111111100100100100011;    //sigmoid(11.937500) ≈ 0.999993
			8'b11000000: sigmoid_out <= 32'b01111111111111111100110001110101;    //sigmoid(12.000000) ≈ 0.999994
			8'b11000001: sigmoid_out <= 32'b01111111111111111100111110010101;    //sigmoid(12.062500) ≈ 0.999994
			8'b11000010: sigmoid_out <= 32'b01111111111111111101001010000100;    //sigmoid(12.125000) ≈ 0.999995
			8'b11000011: sigmoid_out <= 32'b01111111111111111101010101000101;    //sigmoid(12.187500) ≈ 0.999995
			8'b11000100: sigmoid_out <= 32'b01111111111111111101011111011100;    //sigmoid(12.250000) ≈ 0.999995
			8'b11000101: sigmoid_out <= 32'b01111111111111111101101001001011;    //sigmoid(12.312500) ≈ 0.999996
			8'b11000110: sigmoid_out <= 32'b01111111111111111101110010010100;    //sigmoid(12.375000) ≈ 0.999996
			8'b11000111: sigmoid_out <= 32'b01111111111111111101111010111001;    //sigmoid(12.437500) ≈ 0.999996
			8'b11001000: sigmoid_out <= 32'b01111111111111111110000010111101;    //sigmoid(12.500000) ≈ 0.999996
			8'b11001001: sigmoid_out <= 32'b01111111111111111110001010100010;    //sigmoid(12.562500) ≈ 0.999996
			8'b11001010: sigmoid_out <= 32'b01111111111111111110010001101001;    //sigmoid(12.625000) ≈ 0.999997
			8'b11001011: sigmoid_out <= 32'b01111111111111111110011000010101;    //sigmoid(12.687500) ≈ 0.999997
			8'b11001100: sigmoid_out <= 32'b01111111111111111110011110100111;    //sigmoid(12.750000) ≈ 0.999997
			8'b11001101: sigmoid_out <= 32'b01111111111111111110100100100001;    //sigmoid(12.812500) ≈ 0.999997
			8'b11001110: sigmoid_out <= 32'b01111111111111111110101010000100;    //sigmoid(12.875000) ≈ 0.999997
			8'b11001111: sigmoid_out <= 32'b01111111111111111110101111010001;    //sigmoid(12.937500) ≈ 0.999998
			8'b11010000: sigmoid_out <= 32'b01111111111111111110110100001010;    //sigmoid(13.000000) ≈ 0.999998
			8'b11010001: sigmoid_out <= 32'b01111111111111111110111000110000;    //sigmoid(13.062500) ≈ 0.999998
			8'b11010010: sigmoid_out <= 32'b01111111111111111110111101000100;    //sigmoid(13.125000) ≈ 0.999998
			8'b11010011: sigmoid_out <= 32'b01111111111111111111000001001000;    //sigmoid(13.187500) ≈ 0.999998
			8'b11010100: sigmoid_out <= 32'b01111111111111111111000100111100;    //sigmoid(13.250000) ≈ 0.999998
			8'b11010101: sigmoid_out <= 32'b01111111111111111111001000100001;    //sigmoid(13.312500) ≈ 0.999998
			8'b11010110: sigmoid_out <= 32'b01111111111111111111001011111000;    //sigmoid(13.375000) ≈ 0.999998
			8'b11010111: sigmoid_out <= 32'b01111111111111111111001111000010;    //sigmoid(13.437500) ≈ 0.999999
			8'b11011000: sigmoid_out <= 32'b01111111111111111111010010000000;    //sigmoid(13.500000) ≈ 0.999999
			8'b11011001: sigmoid_out <= 32'b01111111111111111111010100110010;    //sigmoid(13.562500) ≈ 0.999999
			8'b11011010: sigmoid_out <= 32'b01111111111111111111010111011010;    //sigmoid(13.625000) ≈ 0.999999
			8'b11011011: sigmoid_out <= 32'b01111111111111111111011001110111;    //sigmoid(13.687500) ≈ 0.999999
			8'b11011100: sigmoid_out <= 32'b01111111111111111111011100001011;    //sigmoid(13.750000) ≈ 0.999999
			8'b11011101: sigmoid_out <= 32'b01111111111111111111011110010110;    //sigmoid(13.812500) ≈ 0.999999
			8'b11011110: sigmoid_out <= 32'b01111111111111111111100000011001;    //sigmoid(13.875000) ≈ 0.999999
			8'b11011111: sigmoid_out <= 32'b01111111111111111111100010010011;    //sigmoid(13.937500) ≈ 0.999999
			8'b11100000: sigmoid_out <= 32'b01111111111111111111100100000110;    //sigmoid(14.000000) ≈ 0.999999
			8'b11100001: sigmoid_out <= 32'b01111111111111111111100101110010;    //sigmoid(14.062500) ≈ 0.999999
			8'b11100010: sigmoid_out <= 32'b01111111111111111111100111011000;    //sigmoid(14.125000) ≈ 0.999999
			8'b11100011: sigmoid_out <= 32'b01111111111111111111101000111000;    //sigmoid(14.187500) ≈ 0.999999
			8'b11100100: sigmoid_out <= 32'b01111111111111111111101010010001;    //sigmoid(14.250000) ≈ 0.999999
			8'b11100101: sigmoid_out <= 32'b01111111111111111111101011100110;    //sigmoid(14.312500) ≈ 0.999999
			8'b11100110: sigmoid_out <= 32'b01111111111111111111101100110101;    //sigmoid(14.375000) ≈ 0.999999
			8'b11100111: sigmoid_out <= 32'b01111111111111111111101101111111;    //sigmoid(14.437500) ≈ 0.999999
			8'b11101000: sigmoid_out <= 32'b01111111111111111111101111000101;    //sigmoid(14.500000) ≈ 0.999999
			8'b11101001: sigmoid_out <= 32'b01111111111111111111110000000111;    //sigmoid(14.562500) ≈ 1.000000
			8'b11101010: sigmoid_out <= 32'b01111111111111111111110001000100;    //sigmoid(14.625000) ≈ 1.000000
			8'b11101011: sigmoid_out <= 32'b01111111111111111111110001111110;    //sigmoid(14.687500) ≈ 1.000000
			8'b11101100: sigmoid_out <= 32'b01111111111111111111110010110100;    //sigmoid(14.750000) ≈ 1.000000
			8'b11101101: sigmoid_out <= 32'b01111111111111111111110011101000;    //sigmoid(14.812500) ≈ 1.000000
			8'b11101110: sigmoid_out <= 32'b01111111111111111111110100011000;    //sigmoid(14.875000) ≈ 1.000000
			8'b11101111: sigmoid_out <= 32'b01111111111111111111110101000101;    //sigmoid(14.937500) ≈ 1.000000
			8'b11110000: sigmoid_out <= 32'b01111111111111111111110101101111;    //sigmoid(15.000000) ≈ 1.000000
			8'b11110001: sigmoid_out <= 32'b01111111111111111111110110010111;    //sigmoid(15.062500) ≈ 1.000000
			8'b11110010: sigmoid_out <= 32'b01111111111111111111110110111100;    //sigmoid(15.125000) ≈ 1.000000
			8'b11110011: sigmoid_out <= 32'b01111111111111111111110111011111;    //sigmoid(15.187500) ≈ 1.000000
			8'b11110100: sigmoid_out <= 32'b01111111111111111111111000000000;    //sigmoid(15.250000) ≈ 1.000000
			8'b11110101: sigmoid_out <= 32'b01111111111111111111111000011111;    //sigmoid(15.312500) ≈ 1.000000
			8'b11110110: sigmoid_out <= 32'b01111111111111111111111000111101;    //sigmoid(15.375000) ≈ 1.000000
			8'b11110111: sigmoid_out <= 32'b01111111111111111111111001011000;    //sigmoid(15.437500) ≈ 1.000000
			8'b11111000: sigmoid_out <= 32'b01111111111111111111111001110010;    //sigmoid(15.500000) ≈ 1.000000
			8'b11111001: sigmoid_out <= 32'b01111111111111111111111010001010;    //sigmoid(15.562500) ≈ 1.000000
			8'b11111010: sigmoid_out <= 32'b01111111111111111111111010100000;    //sigmoid(15.625000) ≈ 1.000000
			8'b11111011: sigmoid_out <= 32'b01111111111111111111111010110110;    //sigmoid(15.687500) ≈ 1.000000
			8'b11111100: sigmoid_out <= 32'b01111111111111111111111011001010;    //sigmoid(15.750000) ≈ 1.000000
			8'b11111101: sigmoid_out <= 32'b01111111111111111111111011011100;    //sigmoid(15.812500) ≈ 1.000000
			8'b11111110: sigmoid_out <= 32'b01111111111111111111111011101110;    //sigmoid(15.875000) ≈ 1.000000
			8'b11111111: sigmoid_out <= 32'b01111111111111111111111011111111;    //sigmoid(15.937500) ≈ 1.000000

        endcase
    end
endmodule