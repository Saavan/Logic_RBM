//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
//
// Create Date: 2019-07-08 15:58:18.364777
// Design Name: vanilla
// Module Name: sigmoidLUT_in8b4p_out6b5p
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 8 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
//
// Additional Comments: Generated by LUT_generator_sigmoid.py
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_in8b4p_out6b5p #(
    parameter PRECISION_INPUT_BITS = 8,
    parameter PRECISION_OUTPUT_BITS = 6
)(
    input[PRECISION_INPUT_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_OUTPUT_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			8'b00000000: sigmoid_out <= 6'b010000;    //sigmoid(0.000000) ≈ 0.500000
			8'b00000001: sigmoid_out <= 6'b010000;    //sigmoid(0.062500) ≈ 0.500000
			8'b00000010: sigmoid_out <= 6'b010001;    //sigmoid(0.125000) ≈ 0.531250
			8'b00000011: sigmoid_out <= 6'b010001;    //sigmoid(0.187500) ≈ 0.531250
			8'b00000100: sigmoid_out <= 6'b010010;    //sigmoid(0.250000) ≈ 0.562500
			8'b00000101: sigmoid_out <= 6'b010010;    //sigmoid(0.312500) ≈ 0.562500
			8'b00000110: sigmoid_out <= 6'b010011;    //sigmoid(0.375000) ≈ 0.593750
			8'b00000111: sigmoid_out <= 6'b010011;    //sigmoid(0.437500) ≈ 0.593750
			8'b00001000: sigmoid_out <= 6'b010100;    //sigmoid(0.500000) ≈ 0.625000
			8'b00001001: sigmoid_out <= 6'b010100;    //sigmoid(0.562500) ≈ 0.625000
			8'b00001010: sigmoid_out <= 6'b010101;    //sigmoid(0.625000) ≈ 0.656250
			8'b00001011: sigmoid_out <= 6'b010101;    //sigmoid(0.687500) ≈ 0.656250
			8'b00001100: sigmoid_out <= 6'b010110;    //sigmoid(0.750000) ≈ 0.687500
			8'b00001101: sigmoid_out <= 6'b010110;    //sigmoid(0.812500) ≈ 0.687500
			8'b00001110: sigmoid_out <= 6'b010111;    //sigmoid(0.875000) ≈ 0.718750
			8'b00001111: sigmoid_out <= 6'b010111;    //sigmoid(0.937500) ≈ 0.718750
			8'b00010000: sigmoid_out <= 6'b010111;    //sigmoid(1.000000) ≈ 0.718750
			8'b00010001: sigmoid_out <= 6'b011000;    //sigmoid(1.062500) ≈ 0.750000
			8'b00010010: sigmoid_out <= 6'b011000;    //sigmoid(1.125000) ≈ 0.750000
			8'b00010011: sigmoid_out <= 6'b011001;    //sigmoid(1.187500) ≈ 0.781250
			8'b00010100: sigmoid_out <= 6'b011001;    //sigmoid(1.250000) ≈ 0.781250
			8'b00010101: sigmoid_out <= 6'b011001;    //sigmoid(1.312500) ≈ 0.781250
			8'b00010110: sigmoid_out <= 6'b011010;    //sigmoid(1.375000) ≈ 0.812500
			8'b00010111: sigmoid_out <= 6'b011010;    //sigmoid(1.437500) ≈ 0.812500
			8'b00011000: sigmoid_out <= 6'b011010;    //sigmoid(1.500000) ≈ 0.812500
			8'b00011001: sigmoid_out <= 6'b011010;    //sigmoid(1.562500) ≈ 0.812500
			8'b00011010: sigmoid_out <= 6'b011011;    //sigmoid(1.625000) ≈ 0.843750
			8'b00011011: sigmoid_out <= 6'b011011;    //sigmoid(1.687500) ≈ 0.843750
			8'b00011100: sigmoid_out <= 6'b011011;    //sigmoid(1.750000) ≈ 0.843750
			8'b00011101: sigmoid_out <= 6'b011100;    //sigmoid(1.812500) ≈ 0.875000
			8'b00011110: sigmoid_out <= 6'b011100;    //sigmoid(1.875000) ≈ 0.875000
			8'b00011111: sigmoid_out <= 6'b011100;    //sigmoid(1.937500) ≈ 0.875000
			8'b00100000: sigmoid_out <= 6'b011100;    //sigmoid(2.000000) ≈ 0.875000
			8'b00100001: sigmoid_out <= 6'b011100;    //sigmoid(2.062500) ≈ 0.875000
			8'b00100010: sigmoid_out <= 6'b011101;    //sigmoid(2.125000) ≈ 0.906250
			8'b00100011: sigmoid_out <= 6'b011101;    //sigmoid(2.187500) ≈ 0.906250
			8'b00100100: sigmoid_out <= 6'b011101;    //sigmoid(2.250000) ≈ 0.906250
			8'b00100101: sigmoid_out <= 6'b011101;    //sigmoid(2.312500) ≈ 0.906250
			8'b00100110: sigmoid_out <= 6'b011101;    //sigmoid(2.375000) ≈ 0.906250
			8'b00100111: sigmoid_out <= 6'b011101;    //sigmoid(2.437500) ≈ 0.906250
			8'b00101000: sigmoid_out <= 6'b011110;    //sigmoid(2.500000) ≈ 0.937500
			8'b00101001: sigmoid_out <= 6'b011110;    //sigmoid(2.562500) ≈ 0.937500
			8'b00101010: sigmoid_out <= 6'b011110;    //sigmoid(2.625000) ≈ 0.937500
			8'b00101011: sigmoid_out <= 6'b011110;    //sigmoid(2.687500) ≈ 0.937500
			8'b00101100: sigmoid_out <= 6'b011110;    //sigmoid(2.750000) ≈ 0.937500
			8'b00101101: sigmoid_out <= 6'b011110;    //sigmoid(2.812500) ≈ 0.937500
			8'b00101110: sigmoid_out <= 6'b011110;    //sigmoid(2.875000) ≈ 0.937500
			8'b00101111: sigmoid_out <= 6'b011110;    //sigmoid(2.937500) ≈ 0.937500
			8'b00110000: sigmoid_out <= 6'b011110;    //sigmoid(3.000000) ≈ 0.937500
			8'b00110001: sigmoid_out <= 6'b011111;    //sigmoid(3.062500) ≈ 0.968750
			8'b00110010: sigmoid_out <= 6'b011111;    //sigmoid(3.125000) ≈ 0.968750
			8'b00110011: sigmoid_out <= 6'b011111;    //sigmoid(3.187500) ≈ 0.968750
			8'b00110100: sigmoid_out <= 6'b011111;    //sigmoid(3.250000) ≈ 0.968750
			8'b00110101: sigmoid_out <= 6'b011111;    //sigmoid(3.312500) ≈ 0.968750
			8'b00110110: sigmoid_out <= 6'b011111;    //sigmoid(3.375000) ≈ 0.968750
			8'b00110111: sigmoid_out <= 6'b011111;    //sigmoid(3.437500) ≈ 0.968750
			8'b00111000: sigmoid_out <= 6'b011111;    //sigmoid(3.500000) ≈ 0.968750
			8'b00111001: sigmoid_out <= 6'b011111;    //sigmoid(3.562500) ≈ 0.968750
			8'b00111010: sigmoid_out <= 6'b011111;    //sigmoid(3.625000) ≈ 0.968750
			8'b00111011: sigmoid_out <= 6'b011111;    //sigmoid(3.687500) ≈ 0.968750
			8'b00111100: sigmoid_out <= 6'b011111;    //sigmoid(3.750000) ≈ 0.968750
			8'b00111101: sigmoid_out <= 6'b011111;    //sigmoid(3.812500) ≈ 0.968750
			8'b00111110: sigmoid_out <= 6'b011111;    //sigmoid(3.875000) ≈ 0.968750
			8'b00111111: sigmoid_out <= 6'b011111;    //sigmoid(3.937500) ≈ 0.968750
			8'b01000000: sigmoid_out <= 6'b011111;    //sigmoid(4.000000) ≈ 0.968750
			8'b01000001: sigmoid_out <= 6'b011111;    //sigmoid(4.062500) ≈ 0.968750
			8'b01000010: sigmoid_out <= 6'b011111;    //sigmoid(4.125000) ≈ 0.968750
			8'b01000011: sigmoid_out <= 6'b100000;    //sigmoid(4.187500) ≈ 1.000000
			8'b01000100: sigmoid_out <= 6'b100000;    //sigmoid(4.250000) ≈ 1.000000
			8'b01000101: sigmoid_out <= 6'b100000;    //sigmoid(4.312500) ≈ 1.000000
			8'b01000110: sigmoid_out <= 6'b100000;    //sigmoid(4.375000) ≈ 1.000000
			8'b01000111: sigmoid_out <= 6'b100000;    //sigmoid(4.437500) ≈ 1.000000
			8'b01001000: sigmoid_out <= 6'b100000;    //sigmoid(4.500000) ≈ 1.000000
			8'b01001001: sigmoid_out <= 6'b100000;    //sigmoid(4.562500) ≈ 1.000000
			8'b01001010: sigmoid_out <= 6'b100000;    //sigmoid(4.625000) ≈ 1.000000
			8'b01001011: sigmoid_out <= 6'b100000;    //sigmoid(4.687500) ≈ 1.000000
			8'b01001100: sigmoid_out <= 6'b100000;    //sigmoid(4.750000) ≈ 1.000000
			8'b01001101: sigmoid_out <= 6'b100000;    //sigmoid(4.812500) ≈ 1.000000
			8'b01001110: sigmoid_out <= 6'b100000;    //sigmoid(4.875000) ≈ 1.000000
			8'b01001111: sigmoid_out <= 6'b100000;    //sigmoid(4.937500) ≈ 1.000000
			8'b01010000: sigmoid_out <= 6'b100000;    //sigmoid(5.000000) ≈ 1.000000
			8'b01010001: sigmoid_out <= 6'b100000;    //sigmoid(5.062500) ≈ 1.000000
			8'b01010010: sigmoid_out <= 6'b100000;    //sigmoid(5.125000) ≈ 1.000000
			8'b01010011: sigmoid_out <= 6'b100000;    //sigmoid(5.187500) ≈ 1.000000
			8'b01010100: sigmoid_out <= 6'b100000;    //sigmoid(5.250000) ≈ 1.000000
			8'b01010101: sigmoid_out <= 6'b100000;    //sigmoid(5.312500) ≈ 1.000000
			8'b01010110: sigmoid_out <= 6'b100000;    //sigmoid(5.375000) ≈ 1.000000
			8'b01010111: sigmoid_out <= 6'b100000;    //sigmoid(5.437500) ≈ 1.000000
			8'b01011000: sigmoid_out <= 6'b100000;    //sigmoid(5.500000) ≈ 1.000000
			8'b01011001: sigmoid_out <= 6'b100000;    //sigmoid(5.562500) ≈ 1.000000
			8'b01011010: sigmoid_out <= 6'b100000;    //sigmoid(5.625000) ≈ 1.000000
			8'b01011011: sigmoid_out <= 6'b100000;    //sigmoid(5.687500) ≈ 1.000000
			8'b01011100: sigmoid_out <= 6'b100000;    //sigmoid(5.750000) ≈ 1.000000
			8'b01011101: sigmoid_out <= 6'b100000;    //sigmoid(5.812500) ≈ 1.000000
			8'b01011110: sigmoid_out <= 6'b100000;    //sigmoid(5.875000) ≈ 1.000000
			8'b01011111: sigmoid_out <= 6'b100000;    //sigmoid(5.937500) ≈ 1.000000
			8'b01100000: sigmoid_out <= 6'b100000;    //sigmoid(6.000000) ≈ 1.000000
			8'b01100001: sigmoid_out <= 6'b100000;    //sigmoid(6.062500) ≈ 1.000000
			8'b01100010: sigmoid_out <= 6'b100000;    //sigmoid(6.125000) ≈ 1.000000
			8'b01100011: sigmoid_out <= 6'b100000;    //sigmoid(6.187500) ≈ 1.000000
			8'b01100100: sigmoid_out <= 6'b100000;    //sigmoid(6.250000) ≈ 1.000000
			8'b01100101: sigmoid_out <= 6'b100000;    //sigmoid(6.312500) ≈ 1.000000
			8'b01100110: sigmoid_out <= 6'b100000;    //sigmoid(6.375000) ≈ 1.000000
			8'b01100111: sigmoid_out <= 6'b100000;    //sigmoid(6.437500) ≈ 1.000000
			8'b01101000: sigmoid_out <= 6'b100000;    //sigmoid(6.500000) ≈ 1.000000
			8'b01101001: sigmoid_out <= 6'b100000;    //sigmoid(6.562500) ≈ 1.000000
			8'b01101010: sigmoid_out <= 6'b100000;    //sigmoid(6.625000) ≈ 1.000000
			8'b01101011: sigmoid_out <= 6'b100000;    //sigmoid(6.687500) ≈ 1.000000
			8'b01101100: sigmoid_out <= 6'b100000;    //sigmoid(6.750000) ≈ 1.000000
			8'b01101101: sigmoid_out <= 6'b100000;    //sigmoid(6.812500) ≈ 1.000000
			8'b01101110: sigmoid_out <= 6'b100000;    //sigmoid(6.875000) ≈ 1.000000
			8'b01101111: sigmoid_out <= 6'b100000;    //sigmoid(6.937500) ≈ 1.000000
			8'b01110000: sigmoid_out <= 6'b100000;    //sigmoid(7.000000) ≈ 1.000000
			8'b01110001: sigmoid_out <= 6'b100000;    //sigmoid(7.062500) ≈ 1.000000
			8'b01110010: sigmoid_out <= 6'b100000;    //sigmoid(7.125000) ≈ 1.000000
			8'b01110011: sigmoid_out <= 6'b100000;    //sigmoid(7.187500) ≈ 1.000000
			8'b01110100: sigmoid_out <= 6'b100000;    //sigmoid(7.250000) ≈ 1.000000
			8'b01110101: sigmoid_out <= 6'b100000;    //sigmoid(7.312500) ≈ 1.000000
			8'b01110110: sigmoid_out <= 6'b100000;    //sigmoid(7.375000) ≈ 1.000000
			8'b01110111: sigmoid_out <= 6'b100000;    //sigmoid(7.437500) ≈ 1.000000
			8'b01111000: sigmoid_out <= 6'b100000;    //sigmoid(7.500000) ≈ 1.000000
			8'b01111001: sigmoid_out <= 6'b100000;    //sigmoid(7.562500) ≈ 1.000000
			8'b01111010: sigmoid_out <= 6'b100000;    //sigmoid(7.625000) ≈ 1.000000
			8'b01111011: sigmoid_out <= 6'b100000;    //sigmoid(7.687500) ≈ 1.000000
			8'b01111100: sigmoid_out <= 6'b100000;    //sigmoid(7.750000) ≈ 1.000000
			8'b01111101: sigmoid_out <= 6'b100000;    //sigmoid(7.812500) ≈ 1.000000
			8'b01111110: sigmoid_out <= 6'b100000;    //sigmoid(7.875000) ≈ 1.000000
			8'b01111111: sigmoid_out <= 6'b100000;    //sigmoid(7.937500) ≈ 1.000000
			8'b10000000: sigmoid_out <= 6'b100000;    //sigmoid(8.000000) ≈ 1.000000
			8'b10000001: sigmoid_out <= 6'b100000;    //sigmoid(8.062500) ≈ 1.000000
			8'b10000010: sigmoid_out <= 6'b100000;    //sigmoid(8.125000) ≈ 1.000000
			8'b10000011: sigmoid_out <= 6'b100000;    //sigmoid(8.187500) ≈ 1.000000
			8'b10000100: sigmoid_out <= 6'b100000;    //sigmoid(8.250000) ≈ 1.000000
			8'b10000101: sigmoid_out <= 6'b100000;    //sigmoid(8.312500) ≈ 1.000000
			8'b10000110: sigmoid_out <= 6'b100000;    //sigmoid(8.375000) ≈ 1.000000
			8'b10000111: sigmoid_out <= 6'b100000;    //sigmoid(8.437500) ≈ 1.000000
			8'b10001000: sigmoid_out <= 6'b100000;    //sigmoid(8.500000) ≈ 1.000000
			8'b10001001: sigmoid_out <= 6'b100000;    //sigmoid(8.562500) ≈ 1.000000
			8'b10001010: sigmoid_out <= 6'b100000;    //sigmoid(8.625000) ≈ 1.000000
			8'b10001011: sigmoid_out <= 6'b100000;    //sigmoid(8.687500) ≈ 1.000000
			8'b10001100: sigmoid_out <= 6'b100000;    //sigmoid(8.750000) ≈ 1.000000
			8'b10001101: sigmoid_out <= 6'b100000;    //sigmoid(8.812500) ≈ 1.000000
			8'b10001110: sigmoid_out <= 6'b100000;    //sigmoid(8.875000) ≈ 1.000000
			8'b10001111: sigmoid_out <= 6'b100000;    //sigmoid(8.937500) ≈ 1.000000
			8'b10010000: sigmoid_out <= 6'b100000;    //sigmoid(9.000000) ≈ 1.000000
			8'b10010001: sigmoid_out <= 6'b100000;    //sigmoid(9.062500) ≈ 1.000000
			8'b10010010: sigmoid_out <= 6'b100000;    //sigmoid(9.125000) ≈ 1.000000
			8'b10010011: sigmoid_out <= 6'b100000;    //sigmoid(9.187500) ≈ 1.000000
			8'b10010100: sigmoid_out <= 6'b100000;    //sigmoid(9.250000) ≈ 1.000000
			8'b10010101: sigmoid_out <= 6'b100000;    //sigmoid(9.312500) ≈ 1.000000
			8'b10010110: sigmoid_out <= 6'b100000;    //sigmoid(9.375000) ≈ 1.000000
			8'b10010111: sigmoid_out <= 6'b100000;    //sigmoid(9.437500) ≈ 1.000000
			8'b10011000: sigmoid_out <= 6'b100000;    //sigmoid(9.500000) ≈ 1.000000
			8'b10011001: sigmoid_out <= 6'b100000;    //sigmoid(9.562500) ≈ 1.000000
			8'b10011010: sigmoid_out <= 6'b100000;    //sigmoid(9.625000) ≈ 1.000000
			8'b10011011: sigmoid_out <= 6'b100000;    //sigmoid(9.687500) ≈ 1.000000
			8'b10011100: sigmoid_out <= 6'b100000;    //sigmoid(9.750000) ≈ 1.000000
			8'b10011101: sigmoid_out <= 6'b100000;    //sigmoid(9.812500) ≈ 1.000000
			8'b10011110: sigmoid_out <= 6'b100000;    //sigmoid(9.875000) ≈ 1.000000
			8'b10011111: sigmoid_out <= 6'b100000;    //sigmoid(9.937500) ≈ 1.000000
			8'b10100000: sigmoid_out <= 6'b100000;    //sigmoid(10.000000) ≈ 1.000000
			8'b10100001: sigmoid_out <= 6'b100000;    //sigmoid(10.062500) ≈ 1.000000
			8'b10100010: sigmoid_out <= 6'b100000;    //sigmoid(10.125000) ≈ 1.000000
			8'b10100011: sigmoid_out <= 6'b100000;    //sigmoid(10.187500) ≈ 1.000000
			8'b10100100: sigmoid_out <= 6'b100000;    //sigmoid(10.250000) ≈ 1.000000
			8'b10100101: sigmoid_out <= 6'b100000;    //sigmoid(10.312500) ≈ 1.000000
			8'b10100110: sigmoid_out <= 6'b100000;    //sigmoid(10.375000) ≈ 1.000000
			8'b10100111: sigmoid_out <= 6'b100000;    //sigmoid(10.437500) ≈ 1.000000
			8'b10101000: sigmoid_out <= 6'b100000;    //sigmoid(10.500000) ≈ 1.000000
			8'b10101001: sigmoid_out <= 6'b100000;    //sigmoid(10.562500) ≈ 1.000000
			8'b10101010: sigmoid_out <= 6'b100000;    //sigmoid(10.625000) ≈ 1.000000
			8'b10101011: sigmoid_out <= 6'b100000;    //sigmoid(10.687500) ≈ 1.000000
			8'b10101100: sigmoid_out <= 6'b100000;    //sigmoid(10.750000) ≈ 1.000000
			8'b10101101: sigmoid_out <= 6'b100000;    //sigmoid(10.812500) ≈ 1.000000
			8'b10101110: sigmoid_out <= 6'b100000;    //sigmoid(10.875000) ≈ 1.000000
			8'b10101111: sigmoid_out <= 6'b100000;    //sigmoid(10.937500) ≈ 1.000000
			8'b10110000: sigmoid_out <= 6'b100000;    //sigmoid(11.000000) ≈ 1.000000
			8'b10110001: sigmoid_out <= 6'b100000;    //sigmoid(11.062500) ≈ 1.000000
			8'b10110010: sigmoid_out <= 6'b100000;    //sigmoid(11.125000) ≈ 1.000000
			8'b10110011: sigmoid_out <= 6'b100000;    //sigmoid(11.187500) ≈ 1.000000
			8'b10110100: sigmoid_out <= 6'b100000;    //sigmoid(11.250000) ≈ 1.000000
			8'b10110101: sigmoid_out <= 6'b100000;    //sigmoid(11.312500) ≈ 1.000000
			8'b10110110: sigmoid_out <= 6'b100000;    //sigmoid(11.375000) ≈ 1.000000
			8'b10110111: sigmoid_out <= 6'b100000;    //sigmoid(11.437500) ≈ 1.000000
			8'b10111000: sigmoid_out <= 6'b100000;    //sigmoid(11.500000) ≈ 1.000000
			8'b10111001: sigmoid_out <= 6'b100000;    //sigmoid(11.562500) ≈ 1.000000
			8'b10111010: sigmoid_out <= 6'b100000;    //sigmoid(11.625000) ≈ 1.000000
			8'b10111011: sigmoid_out <= 6'b100000;    //sigmoid(11.687500) ≈ 1.000000
			8'b10111100: sigmoid_out <= 6'b100000;    //sigmoid(11.750000) ≈ 1.000000
			8'b10111101: sigmoid_out <= 6'b100000;    //sigmoid(11.812500) ≈ 1.000000
			8'b10111110: sigmoid_out <= 6'b100000;    //sigmoid(11.875000) ≈ 1.000000
			8'b10111111: sigmoid_out <= 6'b100000;    //sigmoid(11.937500) ≈ 1.000000
			8'b11000000: sigmoid_out <= 6'b100000;    //sigmoid(12.000000) ≈ 1.000000
			8'b11000001: sigmoid_out <= 6'b100000;    //sigmoid(12.062500) ≈ 1.000000
			8'b11000010: sigmoid_out <= 6'b100000;    //sigmoid(12.125000) ≈ 1.000000
			8'b11000011: sigmoid_out <= 6'b100000;    //sigmoid(12.187500) ≈ 1.000000
			8'b11000100: sigmoid_out <= 6'b100000;    //sigmoid(12.250000) ≈ 1.000000
			8'b11000101: sigmoid_out <= 6'b100000;    //sigmoid(12.312500) ≈ 1.000000
			8'b11000110: sigmoid_out <= 6'b100000;    //sigmoid(12.375000) ≈ 1.000000
			8'b11000111: sigmoid_out <= 6'b100000;    //sigmoid(12.437500) ≈ 1.000000
			8'b11001000: sigmoid_out <= 6'b100000;    //sigmoid(12.500000) ≈ 1.000000
			8'b11001001: sigmoid_out <= 6'b100000;    //sigmoid(12.562500) ≈ 1.000000
			8'b11001010: sigmoid_out <= 6'b100000;    //sigmoid(12.625000) ≈ 1.000000
			8'b11001011: sigmoid_out <= 6'b100000;    //sigmoid(12.687500) ≈ 1.000000
			8'b11001100: sigmoid_out <= 6'b100000;    //sigmoid(12.750000) ≈ 1.000000
			8'b11001101: sigmoid_out <= 6'b100000;    //sigmoid(12.812500) ≈ 1.000000
			8'b11001110: sigmoid_out <= 6'b100000;    //sigmoid(12.875000) ≈ 1.000000
			8'b11001111: sigmoid_out <= 6'b100000;    //sigmoid(12.937500) ≈ 1.000000
			8'b11010000: sigmoid_out <= 6'b100000;    //sigmoid(13.000000) ≈ 1.000000
			8'b11010001: sigmoid_out <= 6'b100000;    //sigmoid(13.062500) ≈ 1.000000
			8'b11010010: sigmoid_out <= 6'b100000;    //sigmoid(13.125000) ≈ 1.000000
			8'b11010011: sigmoid_out <= 6'b100000;    //sigmoid(13.187500) ≈ 1.000000
			8'b11010100: sigmoid_out <= 6'b100000;    //sigmoid(13.250000) ≈ 1.000000
			8'b11010101: sigmoid_out <= 6'b100000;    //sigmoid(13.312500) ≈ 1.000000
			8'b11010110: sigmoid_out <= 6'b100000;    //sigmoid(13.375000) ≈ 1.000000
			8'b11010111: sigmoid_out <= 6'b100000;    //sigmoid(13.437500) ≈ 1.000000
			8'b11011000: sigmoid_out <= 6'b100000;    //sigmoid(13.500000) ≈ 1.000000
			8'b11011001: sigmoid_out <= 6'b100000;    //sigmoid(13.562500) ≈ 1.000000
			8'b11011010: sigmoid_out <= 6'b100000;    //sigmoid(13.625000) ≈ 1.000000
			8'b11011011: sigmoid_out <= 6'b100000;    //sigmoid(13.687500) ≈ 1.000000
			8'b11011100: sigmoid_out <= 6'b100000;    //sigmoid(13.750000) ≈ 1.000000
			8'b11011101: sigmoid_out <= 6'b100000;    //sigmoid(13.812500) ≈ 1.000000
			8'b11011110: sigmoid_out <= 6'b100000;    //sigmoid(13.875000) ≈ 1.000000
			8'b11011111: sigmoid_out <= 6'b100000;    //sigmoid(13.937500) ≈ 1.000000
			8'b11100000: sigmoid_out <= 6'b100000;    //sigmoid(14.000000) ≈ 1.000000
			8'b11100001: sigmoid_out <= 6'b100000;    //sigmoid(14.062500) ≈ 1.000000
			8'b11100010: sigmoid_out <= 6'b100000;    //sigmoid(14.125000) ≈ 1.000000
			8'b11100011: sigmoid_out <= 6'b100000;    //sigmoid(14.187500) ≈ 1.000000
			8'b11100100: sigmoid_out <= 6'b100000;    //sigmoid(14.250000) ≈ 1.000000
			8'b11100101: sigmoid_out <= 6'b100000;    //sigmoid(14.312500) ≈ 1.000000
			8'b11100110: sigmoid_out <= 6'b100000;    //sigmoid(14.375000) ≈ 1.000000
			8'b11100111: sigmoid_out <= 6'b100000;    //sigmoid(14.437500) ≈ 1.000000
			8'b11101000: sigmoid_out <= 6'b100000;    //sigmoid(14.500000) ≈ 1.000000
			8'b11101001: sigmoid_out <= 6'b100000;    //sigmoid(14.562500) ≈ 1.000000
			8'b11101010: sigmoid_out <= 6'b100000;    //sigmoid(14.625000) ≈ 1.000000
			8'b11101011: sigmoid_out <= 6'b100000;    //sigmoid(14.687500) ≈ 1.000000
			8'b11101100: sigmoid_out <= 6'b100000;    //sigmoid(14.750000) ≈ 1.000000
			8'b11101101: sigmoid_out <= 6'b100000;    //sigmoid(14.812500) ≈ 1.000000
			8'b11101110: sigmoid_out <= 6'b100000;    //sigmoid(14.875000) ≈ 1.000000
			8'b11101111: sigmoid_out <= 6'b100000;    //sigmoid(14.937500) ≈ 1.000000
			8'b11110000: sigmoid_out <= 6'b100000;    //sigmoid(15.000000) ≈ 1.000000
			8'b11110001: sigmoid_out <= 6'b100000;    //sigmoid(15.062500) ≈ 1.000000
			8'b11110010: sigmoid_out <= 6'b100000;    //sigmoid(15.125000) ≈ 1.000000
			8'b11110011: sigmoid_out <= 6'b100000;    //sigmoid(15.187500) ≈ 1.000000
			8'b11110100: sigmoid_out <= 6'b100000;    //sigmoid(15.250000) ≈ 1.000000
			8'b11110101: sigmoid_out <= 6'b100000;    //sigmoid(15.312500) ≈ 1.000000
			8'b11110110: sigmoid_out <= 6'b100000;    //sigmoid(15.375000) ≈ 1.000000
			8'b11110111: sigmoid_out <= 6'b100000;    //sigmoid(15.437500) ≈ 1.000000
			8'b11111000: sigmoid_out <= 6'b100000;    //sigmoid(15.500000) ≈ 1.000000
			8'b11111001: sigmoid_out <= 6'b100000;    //sigmoid(15.562500) ≈ 1.000000
			8'b11111010: sigmoid_out <= 6'b100000;    //sigmoid(15.625000) ≈ 1.000000
			8'b11111011: sigmoid_out <= 6'b100000;    //sigmoid(15.687500) ≈ 1.000000
			8'b11111100: sigmoid_out <= 6'b100000;    //sigmoid(15.750000) ≈ 1.000000
			8'b11111101: sigmoid_out <= 6'b100000;    //sigmoid(15.812500) ≈ 1.000000
			8'b11111110: sigmoid_out <= 6'b100000;    //sigmoid(15.875000) ≈ 1.000000
			8'b11111111: sigmoid_out <= 6'b100000;    //sigmoid(15.937500) ≈ 1.000000

        endcase
    end
endmodule