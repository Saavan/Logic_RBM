//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
//
// Create Date: 2019-07-08 11:13:08.772110
// Design Name: vanilla
// Module Name: sigmoidLUT_in8b4p_out64b63p
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 8 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
//
// Additional Comments: Generated by LUT_generator_sigmoid.py
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_in8b4p_out64b63p #(
    parameter PRECISION_INPUT_BITS = 8,
    parameter PRECISION_OUTPUT_BITS = 64
)(
    input[PRECISION_INPUT_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_OUTPUT_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			8'b00000000: sigmoid_out <= 64'b0100000000000000000000000000000000000000000000000000000000000000;    //sigmoid(0.000000) ≈ 0.500000
			8'b00000001: sigmoid_out <= 64'b0100000111111111110101010101100110011001001010110001110000000000;    //sigmoid(0.062500) ≈ 0.515620
			8'b00000010: sigmoid_out <= 64'b0100001111111110101010110011001011111100000001100001110000000000;    //sigmoid(0.125000) ≈ 0.531209
			8'b00000011: sigmoid_out <= 64'b0100010111111011100001000000100100011111111011000010010000000000;    //sigmoid(0.187500) ≈ 0.546738
			8'b00000100: sigmoid_out <= 64'b0100011111110101011001100100101011110001001011100000110000000000;    //sigmoid(0.250000) ≈ 0.562177
			8'b00000101: sigmoid_out <= 64'b0100100111101011010111100011110110001000010001100001010000000000;    //sigmoid(0.312500) ≈ 0.577495
			8'b00000110: sigmoid_out <= 64'b0100101111011100011111111100100000011101111110111011100000000000;    //sigmoid(0.375000) ≈ 0.592667
			8'b00000111: sigmoid_out <= 64'b0100110111000111111010000010000010110101001111100100110000000000;    //sigmoid(0.437500) ≈ 0.607663
			8'b00001000: sigmoid_out <= 64'b0100111110101100101111110101001101001101000011100100010000000000;    //sigmoid(0.500000) ≈ 0.622459
			8'b00001001: sigmoid_out <= 64'b0101000110001010001110011001111001101011010010000100010000000000;    //sigmoid(0.562500) ≈ 0.637031
			8'b00001010: sigmoid_out <= 64'b0101001101011111100110001010000011101010011001010000110000000000;    //sigmoid(0.625000) ≈ 0.651355
			8'b00001011: sigmoid_out <= 64'b0101010100101100001011000101011000011101100001100000100000000000;    //sigmoid(0.687500) ≈ 0.665411
			8'b00001100: sigmoid_out <= 64'b0101011011101111010100111101111010001100100011111011000000000000;    //sigmoid(0.750000) ≈ 0.679179
			8'b00001101: sigmoid_out <= 64'b0101100010101000011111100001010010110011001111000011100000000000;    //sigmoid(0.812500) ≈ 0.692642
			8'b00001110: sigmoid_out <= 64'b0101101001010111001010011110111001001000100000000011100000000000;    //sigmoid(0.875000) ≈ 0.705785
			8'b00001111: sigmoid_out <= 64'b0101101111111010111001101010101110010111001001001101110000000000;    //sigmoid(0.937500) ≈ 0.718594
			8'b00010000: sigmoid_out <= 64'b0101110110010011010100111101011101010110100010101111010000000000;    //sigmoid(1.000000) ≈ 0.731059
			8'b00010001: sigmoid_out <= 64'b0101111100100000001000010001101000110110010001110101110000000000;    //sigmoid(1.062500) ≈ 0.743168
			8'b00010010: sigmoid_out <= 64'b0110000010100001000011011110010111101101101010010110110000000000;    //sigmoid(1.125000) ≈ 0.754915
			8'b00010011: sigmoid_out <= 64'b0110001000010101111010001111110000010111111011000010000000000000;    //sigmoid(1.187500) ≈ 0.766294
			8'b00010100: sigmoid_out <= 64'b0110001101111110100011111101010101110111000111110010100000000000;    //sigmoid(1.250000) ≈ 0.777300
			8'b00010101: sigmoid_out <= 64'b0110010011011010111011011110111001100100011001111001000000000000;    //sigmoid(1.312500) ≈ 0.787931
			8'b00010110: sigmoid_out <= 64'b0110011000101010111110111111110100111110111000101011100000000000;    //sigmoid(1.375000) ≈ 0.798187
			8'b00010111: sigmoid_out <= 64'b0110011101101110101111110001011110010110111010000101110000000000;    //sigmoid(1.437500) ≈ 0.808067
			8'b00011000: sigmoid_out <= 64'b0110100010100110010001111100101010100101111001000101000000000000;    //sigmoid(1.500000) ≈ 0.817574
			8'b00011001: sigmoid_out <= 64'b0110100111010001101100010010101101100000001000011011100000000000;    //sigmoid(1.562500) ≈ 0.826712
			8'b00011010: sigmoid_out <= 64'b0110101011110001000111111110001000011010010100110011010000000000;    //sigmoid(1.625000) ≈ 0.835484
			8'b00011011: sigmoid_out <= 64'b0110110000000100110000010011010101011100111110000100010000000000;    //sigmoid(1.687500) ≈ 0.843895
			8'b00011100: sigmoid_out <= 64'b0110110100001100110010100001011100011000010000000010110000000000;    //sigmoid(1.750000) ≈ 0.851953
			8'b00011101: sigmoid_out <= 64'b0110111000001001011101100011011011111111100101110000000000000000;    //sigmoid(1.812500) ≈ 0.859664
			8'b00011110: sigmoid_out <= 64'b0110111011111011000001110001110001101000000010101111010000000000;    //sigmoid(1.875000) ≈ 0.867036
			8'b00011111: sigmoid_out <= 64'b0110111111100001110000110100100110011011000010001101110000000000;    //sigmoid(1.937500) ≈ 0.874077
			8'b00100000: sigmoid_out <= 64'b0111000010111101111101010110101000101001111001110010010000000000;    //sigmoid(2.000000) ≈ 0.880797
			8'b00100001: sigmoid_out <= 64'b0111000110001111111010111000110101110000000111101101010000000000;    //sigmoid(2.062500) ≈ 0.887205
			8'b00100010: sigmoid_out <= 64'b0111001001010111111101100110111000011011001101101110000000000000;    //sigmoid(2.125000) ≈ 0.893309
			8'b00100011: sigmoid_out <= 64'b0111001100010110011010001100011101000001001000110010100000000000;    //sigmoid(2.187500) ≈ 0.899121
			8'b00100100: sigmoid_out <= 64'b0111001111001011100101101011011101001000100110101101010000000000;    //sigmoid(2.250000) ≈ 0.904651
			8'b00100101: sigmoid_out <= 64'b0111010001110111110101010011000010101010110101110010110000000000;    //sigmoid(2.312500) ≈ 0.909907
			8'b00100110: sigmoid_out <= 64'b0111010100011011011110010111100001100011000100101111010000000000;    //sigmoid(2.375000) ≈ 0.914901
			8'b00100111: sigmoid_out <= 64'b0111010110110110110110001011000110110101101010110000000000000000;    //sigmoid(2.437500) ≈ 0.919643
			8'b00101000: sigmoid_out <= 64'b0111011001001010010001110111011011010110010110111110000000000000;    //sigmoid(2.500000) ≈ 0.924142
			8'b00101001: sigmoid_out <= 64'b0111011011010110000110010111110111011010001001000101100000000000;    //sigmoid(2.562500) ≈ 0.928409
			8'b00101010: sigmoid_out <= 64'b0111011101011010101000010100100101001101000101111000010000000000;    //sigmoid(2.625000) ≈ 0.932453
			8'b00101011: sigmoid_out <= 64'b0111011111011000001011111110001110110110001001000011110000000000;    //sigmoid(2.687500) ≈ 0.936285
			8'b00101100: sigmoid_out <= 64'b0111100001001111000101001010010101001001110010001111000000000000;    //sigmoid(2.750000) ≈ 0.939913
			8'b00101101: sigmoid_out <= 64'b0111100010111111100111010000001100001000000101011111000000000000;    //sigmoid(2.812500) ≈ 0.943348
			8'b00101110: sigmoid_out <= 64'b0111100100101010000101000110011010000001100100010111110000000000;    //sigmoid(2.875000) ≈ 0.946597
			8'b00101111: sigmoid_out <= 64'b0111100110001110110001000000110110000000111000000101000000000000;    //sigmoid(2.937500) ≈ 0.949669
			8'b00110000: sigmoid_out <= 64'b0111100111101101111100101111000011011011111010101111010000000000;    //sigmoid(3.000000) ≈ 0.952574
			8'b00110001: sigmoid_out <= 64'b0111101001000111111001011011000110110110000010001111100000000000;    //sigmoid(3.062500) ≈ 0.955319
			8'b00110010: sigmoid_out <= 64'b0111101010011100110111101000110010000101000011010110000000000000;    //sigmoid(3.125000) ≈ 0.957912
			8'b00110011: sigmoid_out <= 64'b0111101011101101000111010101000100110100011110001000010000000000;    //sigmoid(3.187500) ≈ 0.960361
			8'b00110100: sigmoid_out <= 64'b0111101100111000110111110101111111001100001110001111010000000000;    //sigmoid(3.250000) ≈ 0.962673
			8'b00110101: sigmoid_out <= 64'b0111101110000000010111111010100100001010111101101001000000000000;    //sigmoid(3.312500) ≈ 0.964855
			8'b00110110: sigmoid_out <= 64'b0111101111000011110101101011001001101110101000110001110000000000;    //sigmoid(3.375000) ≈ 0.966914
			8'b00110111: sigmoid_out <= 64'b0111110000000011011110101001110100110000110000110101000000000000;    //sigmoid(3.437500) ≈ 0.968856
			8'b00111000: sigmoid_out <= 64'b0111110000111111011111110010111111000110011010100100110000000000;    //sigmoid(3.500000) ≈ 0.970688
			8'b00111001: sigmoid_out <= 64'b0111110001111000000101011110000101111110000101001011000000000000;    //sigmoid(3.562500) ≈ 0.972415
			8'b00111010: sigmoid_out <= 64'b0111110010101101011011011110011111011111010101111111100000000000;    //sigmoid(3.625000) ≈ 0.974043
			8'b00111011: sigmoid_out <= 64'b0111110011011111101101000100010101111001101001001111100000000000;    //sigmoid(3.687500) ≈ 0.975577
			8'b00111100: sigmoid_out <= 64'b0111110100001111000100111101100111011000000110111011010000000000;    //sigmoid(3.750000) ≈ 0.977023
			8'b00111101: sigmoid_out <= 64'b0111110100111011101101010111001001011000100111000101100000000000;    //sigmoid(3.812500) ≈ 0.978385
			8'b00111110: sigmoid_out <= 64'b0111110101100101101111111101101110101011110110010010010000000000;    //sigmoid(3.875000) ≈ 0.979668
			8'b00111111: sigmoid_out <= 64'b0111110110001101010101111111001111001011001100001110110000000000;    //sigmoid(3.937500) ≈ 0.980876
			8'b01000000: sigmoid_out <= 64'b0111110110110010101000001011110000110111100001111010100000000000;    //sigmoid(4.000000) ≈ 0.982014
			8'b01000001: sigmoid_out <= 64'b0111110111010101101110110110110001011010001101001011000000000000;    //sigmoid(4.062500) ≈ 0.983085
			8'b01000010: sigmoid_out <= 64'b0111110111110110110001111000001111100110011100110011000000000000;    //sigmoid(4.125000) ≈ 0.984094
			8'b01000011: sigmoid_out <= 64'b0111111000010101111000101101110100011110100101101110110000000000;    //sigmoid(4.187500) ≈ 0.985043
			8'b01000100: sigmoid_out <= 64'b0111111000110011001010011011111011100100100111111000110000000000;    //sigmoid(4.250000) ≈ 0.985936
			8'b01000101: sigmoid_out <= 64'b0111111001001110101101101110111010000001101010100110000000000000;    //sigmoid(4.312500) ≈ 0.986777
			8'b01000110: sigmoid_out <= 64'b0111111001101000101000111100000100010011001111000100000000000000;    //sigmoid(4.375000) ≈ 0.987568
			8'b01000111: sigmoid_out <= 64'b0111111010000001000010000010110010010000011101010100000000000000;    //sigmoid(4.437500) ≈ 0.988313
			8'b01001000: sigmoid_out <= 64'b0111111010010111111110101101100001011011111110100011110000000000;    //sigmoid(4.500000) ≈ 0.989013
			8'b01001001: sigmoid_out <= 64'b0111111010101101100100010010110101011001110010100100000000000000;    //sigmoid(4.562500) ≈ 0.989672
			8'b01001010: sigmoid_out <= 64'b0111111011000001110111110110010110000010010100001001000000000000;    //sigmoid(4.625000) ≈ 0.990292
			8'b01001011: sigmoid_out <= 64'b0111111011010100111110001001101011101101110111010100000000000000;    //sigmoid(4.687500) ≈ 0.990874
			8'b01001100: sigmoid_out <= 64'b0111111011100110111011101101011001010101010001011011100000000000;    //sigmoid(4.750000) ≈ 0.991423
			8'b01001101: sigmoid_out <= 64'b0111111011110111110100110001110100000101110100010010000000000000;    //sigmoid(4.812500) ≈ 0.991938
			8'b01001110: sigmoid_out <= 64'b0111111100000111101101010111111001000111110000101111000000000000;    //sigmoid(4.875000) ≈ 0.992423
			8'b01001111: sigmoid_out <= 64'b0111111100010110101001010010000000110111110101111101000000000000;    //sigmoid(4.937500) ≈ 0.992879
			8'b01010000: sigmoid_out <= 64'b0111111100100100101100000100110000010100111000111000100000000000;    //sigmoid(5.000000) ≈ 0.993307
			8'b01010001: sigmoid_out <= 64'b0111111100110001111001000111101000000011011101001111000000000000;    //sigmoid(5.062500) ≈ 0.993710
			8'b01010010: sigmoid_out <= 64'b0111111100111110010011100101110001001001111111001101100000000000;    //sigmoid(5.125000) ≈ 0.994089
			8'b01010011: sigmoid_out <= 64'b0111111101001001111110011110101000001000011011111001000000000000;    //sigmoid(5.187500) ≈ 0.994445
			8'b01010100: sigmoid_out <= 64'b0111111101010100111100100110100101101110101111010111110000000000;    //sigmoid(5.250000) ≈ 0.994780
			8'b01010101: sigmoid_out <= 64'b0111111101011111010000100111100101110101110011001100100000000000;    //sigmoid(5.312500) ≈ 0.995095
			8'b01010110: sigmoid_out <= 64'b0111111101101000111101000001101100011110110110100100110000000000;    //sigmoid(5.375000) ≈ 0.995390
			8'b01010111: sigmoid_out <= 64'b0111111101110010000100001011101000111101010100111101000000000000;    //sigmoid(5.437500) ≈ 0.995668
			8'b01011000: sigmoid_out <= 64'b0111111101111010101000010011010111001111010111001000000000000000;    //sigmoid(5.500000) ≈ 0.995930
			8'b01011001: sigmoid_out <= 64'b0111111110000010101011011110011111101001001111011011100000000000;    //sigmoid(5.562500) ≈ 0.996176
			8'b01011010: sigmoid_out <= 64'b0111111110001010001111101010110100111000000011111011010000000000;    //sigmoid(5.625000) ≈ 0.996406
			8'b01011011: sigmoid_out <= 64'b0111111110010001010110101110110000011111111001001000000000000000;    //sigmoid(5.687500) ≈ 0.996623
			8'b01011100: sigmoid_out <= 64'b0111111110011000000010011001101101111001101110001001100000000000;    //sigmoid(5.750000) ≈ 0.996827
			8'b01011101: sigmoid_out <= 64'b0111111110011110010100010100100011110101010111110011010000000000;    //sigmoid(5.812500) ≈ 0.997019
			8'b01011110: sigmoid_out <= 64'b0111111110100100001110000001111100100011100011001010110000000000;    //sigmoid(5.875000) ≈ 0.997199
			8'b01011111: sigmoid_out <= 64'b0111111110101001110000111110101100101100000011001010110000000000;    //sigmoid(5.937500) ≈ 0.997368
			8'b01100000: sigmoid_out <= 64'b0111111110101110111110100010001000110100000101100000010000000000;    //sigmoid(6.000000) ≈ 0.997527
			8'b01100001: sigmoid_out <= 64'b0111111110110011110111111110011001111000100100111010100000000000;    //sigmoid(6.062500) ≈ 0.997677
			8'b01100010: sigmoid_out <= 64'b0111111110111000011110100000110000100000000110100011110000000000;    //sigmoid(6.125000) ≈ 0.997817
			8'b01100011: sigmoid_out <= 64'b0111111110111100110011010001110111001000001000110001110000000000;    //sigmoid(6.187500) ≈ 0.997949
			8'b01100100: sigmoid_out <= 64'b0111111111000000110111010110000011010001000001000010010000000000;    //sigmoid(6.250000) ≈ 0.998073
			8'b01100101: sigmoid_out <= 64'b0111111111000100101011101101100101101011111110110010000000000000;    //sigmoid(6.312500) ≈ 0.998190
			8'b01100110: sigmoid_out <= 64'b0111111111001000010001010100111001101110100000010000000000000000;    //sigmoid(6.375000) ≈ 0.998299
			8'b01100111: sigmoid_out <= 64'b0111111111001011101001000100110011101101111110000010000000000000;    //sigmoid(6.437500) ≈ 0.998402
			8'b01101000: sigmoid_out <= 64'b0111111111001110110011110010101110100110101001110100000000000000;    //sigmoid(6.500000) ≈ 0.998499
			8'b01101001: sigmoid_out <= 64'b0111111111010001110010010000111000110000110100010110000000000000;    //sigmoid(6.562500) ≈ 0.998590
			8'b01101010: sigmoid_out <= 64'b0111111111010100100101001110100000000110100110101110100000000000;    //sigmoid(6.625000) ≈ 0.998675
			8'b01101011: sigmoid_out <= 64'b0111111111010111001101010111111101011101010011000010000000000000;    //sigmoid(6.687500) ≈ 0.998755
			8'b01101100: sigmoid_out <= 64'b0111111111011001101011010110111111010100011000100101000000000000;    //sigmoid(6.750000) ≈ 0.998830
			8'b01101101: sigmoid_out <= 64'b0111111111011011111111110010110011111100110000101010000000000000;    //sigmoid(6.812500) ≈ 0.998901
			8'b01101110: sigmoid_out <= 64'b0111111111011110001011010000010010111010010001001011100000000000;    //sigmoid(6.875000) ≈ 0.998968
			8'b01101111: sigmoid_out <= 64'b0111111111100000001110010010000110000001101011101010010000000000;    //sigmoid(6.937500) ≈ 0.999030
			8'b01110000: sigmoid_out <= 64'b0111111111100010001001011000110001110101001000001111000000000000;    //sigmoid(7.000000) ≈ 0.999089
			8'b01110001: sigmoid_out <= 64'b0111111111100011111101000010111101100000110101101100010000000000;    //sigmoid(7.062500) ≈ 0.999144
			8'b01110010: sigmoid_out <= 64'b0111111111100101101001101101011010011010000001011011010000000000;    //sigmoid(7.125000) ≈ 0.999196
			8'b01110011: sigmoid_out <= 64'b0111111111100111001111110011001011000001100100000011000000000000;    //sigmoid(7.187500) ≈ 0.999245
			8'b01110100: sigmoid_out <= 64'b0111111111101000101111101101101001101100001001100111100000000000;    //sigmoid(7.250000) ≈ 0.999290
			8'b01110101: sigmoid_out <= 64'b0111111111101010001001110100101110110001010111000110000000000000;    //sigmoid(7.312500) ≈ 0.999333
			8'b01110110: sigmoid_out <= 64'b0111111111101011011110011110110110100011001001001000010000000000;    //sigmoid(7.375000) ≈ 0.999374
			8'b01110111: sigmoid_out <= 64'b0111111111101100101110000001000110101111000011100010110000000000;    //sigmoid(7.437500) ≈ 0.999412
			8'b01111000: sigmoid_out <= 64'b0111111111101101111000101111010011101010100011101110010000000000;    //sigmoid(7.500000) ≈ 0.999447
			8'b01111001: sigmoid_out <= 64'b0111111111101110111110111100000101001011100100000100010000000000;    //sigmoid(7.562500) ≈ 0.999481
			8'b01111010: sigmoid_out <= 64'b0111111111110000000000111000111011001110011001110110000000000000;    //sigmoid(7.625000) ≈ 0.999512
			8'b01111011: sigmoid_out <= 64'b0111111111110000111110110110010010001010010010111100100000000000;    //sigmoid(7.687500) ≈ 0.999542
			8'b01111100: sigmoid_out <= 64'b0111111111110001111001000011100110110101010101001100100000000000;    //sigmoid(7.750000) ≈ 0.999569
			8'b01111101: sigmoid_out <= 64'b0111111111110010101111101111011010011000111100111000000000000000;    //sigmoid(7.812500) ≈ 0.999596
			8'b01111110: sigmoid_out <= 64'b0111111111110011100011000111010101110111110100111110010000000000;    //sigmoid(7.875000) ≈ 0.999620
			8'b01111111: sigmoid_out <= 64'b0111111111110100010011011000001101100110000000000011000000000000;    //sigmoid(7.937500) ≈ 0.999643
			8'b10000000: sigmoid_out <= 64'b0111111111110101000000101110000100010100000101101000100000000000;    //sigmoid(8.000000) ≈ 0.999665
			8'b10000001: sigmoid_out <= 64'b0111111111110101101011010100001110001110010101000100010000000000;    //sigmoid(8.062500) ≈ 0.999685
			8'b10000010: sigmoid_out <= 64'b0111111111110110010011010101010011110000001011110100100000000000;    //sigmoid(8.125000) ≈ 0.999704
			8'b10000011: sigmoid_out <= 64'b0111111111110110111000111011010100001101001010101101110000000000;    //sigmoid(8.187500) ≈ 0.999722
			8'b10000100: sigmoid_out <= 64'b0111111111110111011100001111101000001111100010111100000000000000;    //sigmoid(8.250000) ≈ 0.999739
			8'b10000101: sigmoid_out <= 64'b0111111111110111111101011011000100001101100001010101110000000000;    //sigmoid(8.312500) ≈ 0.999755
			8'b10000110: sigmoid_out <= 64'b0111111111111000011100100101111010010101011100011010100000000000;    //sigmoid(8.375000) ≈ 0.999769
			8'b10000111: sigmoid_out <= 64'b0111111111111000111001110111111100110001100110110111100000000000;    //sigmoid(8.437500) ≈ 0.999783
			8'b10001000: sigmoid_out <= 64'b0111111111111001010101011000011111100100000111001100110000000000;    //sigmoid(8.500000) ≈ 0.999797
			8'b10001001: sigmoid_out <= 64'b0111111111111001101111001110011010011011010010011000010000000000;    //sigmoid(8.562500) ≈ 0.999809
			8'b10001010: sigmoid_out <= 64'b0111111111111010000111100000001010011111000110001001110000000000;    //sigmoid(8.625000) ≈ 0.999820
			8'b10001011: sigmoid_out <= 64'b0111111111111010011110010011110011110111111101110101110000000000;    //sigmoid(8.687500) ≈ 0.999831
			8'b10001100: sigmoid_out <= 64'b0111111111111010110011101111000011001111011010110000000000000000;    //sigmoid(8.750000) ≈ 0.999842
			8'b10001101: sigmoid_out <= 64'b0111111111111011000111110111001111001010111000000001000000000000;    //sigmoid(8.812500) ≈ 0.999851
			8'b10001110: sigmoid_out <= 64'b0111111111111011011010110001011001100001000000001100100000000000;    //sigmoid(8.875000) ≈ 0.999860
			8'b10001111: sigmoid_out <= 64'b0111111111111011101100100010010000101001111001100001010000000000;    //sigmoid(8.937500) ≈ 0.999869
			8'b10010000: sigmoid_out <= 64'b0111111111111011111101001110010000101010011100110000010000000000;    //sigmoid(9.000000) ≈ 0.999877
			8'b10010001: sigmoid_out <= 64'b0111111111111100001100111001100100011011001001000010010000000000;    //sigmoid(9.062500) ≈ 0.999884
			8'b10010010: sigmoid_out <= 64'b0111111111111100011011101000000110101010100110010011010000000000;    //sigmoid(9.125000) ≈ 0.999891
			8'b10010011: sigmoid_out <= 64'b0111111111111100101001011101100010111100000110101100010000000000;    //sigmoid(9.187500) ≈ 0.999898
			8'b10010100: sigmoid_out <= 64'b0111111111111100110110011101010110100010010110011011100000000000;    //sigmoid(9.250000) ≈ 0.999904
			8'b10010101: sigmoid_out <= 64'b0111111111111101000010101010110001010110101000101000000000000000;    //sigmoid(9.312500) ≈ 0.999910
			8'b10010110: sigmoid_out <= 64'b0111111111111101001110001000110110101100101110110000100000000000;    //sigmoid(9.375000) ≈ 0.999915
			8'b10010111: sigmoid_out <= 64'b0111111111111101011000111010011110000011100111100111100000000000;    //sigmoid(9.437500) ≈ 0.999920
			8'b10011000: sigmoid_out <= 64'b0111111111111101100011000010010011110011010001110100110000000000;    //sigmoid(9.500000) ≈ 0.999925
			8'b10011001: sigmoid_out <= 64'b0111111111111101101100100010111001110111101101010001110000000000;    //sigmoid(9.562500) ≈ 0.999930
			8'b10011010: sigmoid_out <= 64'b0111111111111101110101011110101000011001010110001011000000000000;    //sigmoid(9.625000) ≈ 0.999934
			8'b10011011: sigmoid_out <= 64'b0111111111111101111101110111101110010011000011101000100000000000;    //sigmoid(9.687500) ≈ 0.999938
			8'b10011100: sigmoid_out <= 64'b0111111111111110000101110000010001110101110011011100110000000000;    //sigmoid(9.750000) ≈ 0.999942
			8'b10011101: sigmoid_out <= 64'b0111111111111110001101001010010001001010001011101100110000000000;    //sigmoid(9.812500) ≈ 0.999945
			8'b10011110: sigmoid_out <= 64'b0111111111111110010100000111100010101111111010101000000000000000;    //sigmoid(9.875000) ≈ 0.999949
			8'b10011111: sigmoid_out <= 64'b0111111111111110011010101001110101111011011100100101110000000000;    //sigmoid(9.937500) ≈ 0.999952
			8'b10100000: sigmoid_out <= 64'b0111111111111110100000110010110011010001101111100010010000000000;    //sigmoid(10.000000) ≈ 0.999955
			8'b10100001: sigmoid_out <= 64'b0111111111111110100110100011111101000010011010101101100000000000;    //sigmoid(10.062500) ≈ 0.999957
			8'b10100010: sigmoid_out <= 64'b0111111111111110101011111110101111100000010001010111000000000000;    //sigmoid(10.125000) ≈ 0.999960
			8'b10100011: sigmoid_out <= 64'b0111111111111110110001000100100001011000010110010010010000000000;    //sigmoid(10.187500) ≈ 0.999962
			8'b10100100: sigmoid_out <= 64'b0111111111111110110101110110100100000111100110001111000000000000;    //sigmoid(10.250000) ≈ 0.999965
			8'b10100101: sigmoid_out <= 64'b0111111111111110111010010110000100001111001110010100110000000000;    //sigmoid(10.312500) ≈ 0.999967
			8'b10100110: sigmoid_out <= 64'b0111111111111110111110100100001001100111110011101000100000000000;    //sigmoid(10.375000) ≈ 0.999969
			8'b10100111: sigmoid_out <= 64'b0111111111111111000010100001110111110011010000110100110000000000;    //sigmoid(10.437500) ≈ 0.999971
			8'b10101000: sigmoid_out <= 64'b0111111111111111000110010000001110001101101110000110010000000000;    //sigmoid(10.500000) ≈ 0.999972
			8'b10101001: sigmoid_out <= 64'b0111111111111111001001110000001000011101010111110110010000000000;    //sigmoid(10.562500) ≈ 0.999974
			8'b10101010: sigmoid_out <= 64'b0111111111111111001101000010011110100001010111110110000000000000;    //sigmoid(10.625000) ≈ 0.999976
			8'b10101011: sigmoid_out <= 64'b0111111111111111010000001000000100111111110100101110100000000000;    //sigmoid(10.687500) ≈ 0.999977
			8'b10101100: sigmoid_out <= 64'b0111111111111111010011000001101101010010111011010101100000000000;    //sigmoid(10.750000) ≈ 0.999979
			8'b10101101: sigmoid_out <= 64'b0111111111111111010101110000000101110101010101000010110000000000;    //sigmoid(10.812500) ≈ 0.999980
			8'b10101110: sigmoid_out <= 64'b0111111111111111011000010011111010001101101110010001110000000000;    //sigmoid(10.875000) ≈ 0.999981
			8'b10101111: sigmoid_out <= 64'b0111111111111111011010101101110011011001110000000011000000000000;    //sigmoid(10.937500) ≈ 0.999982
			8'b10110000: sigmoid_out <= 64'b0111111111111111011100111110010111111000001111010010100000000000;    //sigmoid(11.000000) ≈ 0.999983
			8'b10110001: sigmoid_out <= 64'b0111111111111111011111000110001011110010110100011110010000000000;    //sigmoid(11.062500) ≈ 0.999984
			8'b10110010: sigmoid_out <= 64'b0111111111111111100001000101110001000110111101111111110000000000;    //sigmoid(11.125000) ≈ 0.999985
			8'b10110011: sigmoid_out <= 64'b0111111111111111100010111101100111101110011111011111010000000000;    //sigmoid(11.187500) ≈ 0.999986
			8'b10110100: sigmoid_out <= 64'b0111111111111111100100101110001101100111100000001110100000000000;    //sigmoid(11.250000) ≈ 0.999987
			8'b10110101: sigmoid_out <= 64'b0111111111111111100110010111111110111011111010101101100000000000;    //sigmoid(11.312500) ≈ 0.999988
			8'b10110110: sigmoid_out <= 64'b0111111111111111100111111011010110001000011111000110010000000000;    //sigmoid(11.375000) ≈ 0.999989
			8'b10110111: sigmoid_out <= 64'b0111111111111111101001011000101100000011011010011001010000000000;    //sigmoid(11.437500) ≈ 0.999989
			8'b10111000: sigmoid_out <= 64'b0111111111111111101010110000011000000010100100000100110000000000;    //sigmoid(11.500000) ≈ 0.999990
			8'b10111001: sigmoid_out <= 64'b0111111111111111101100000010110000000001010011100000010000000000;    //sigmoid(11.562500) ≈ 0.999990
			8'b10111010: sigmoid_out <= 64'b0111111111111111101101010000001000100101111110110110010000000000;    //sigmoid(11.625000) ≈ 0.999991
			8'b10111011: sigmoid_out <= 64'b0111111111111111101110011000110101000111000100101100100000000000;    //sigmoid(11.687500) ≈ 0.999992
			8'b10111100: sigmoid_out <= 64'b0111111111111111101111011101000111110000000001101010010000000000;    //sigmoid(11.750000) ≈ 0.999992
			8'b10111101: sigmoid_out <= 64'b0111111111111111110000011101010001100101110011010101010000000000;    //sigmoid(11.812500) ≈ 0.999993
			8'b10111110: sigmoid_out <= 64'b0111111111111111110001011001100010101011001001100001010000000000;    //sigmoid(11.875000) ≈ 0.999993
			8'b10111111: sigmoid_out <= 64'b0111111111111111110010010010001010000100100110111111000000000000;    //sigmoid(11.937500) ≈ 0.999993
			8'b11000000: sigmoid_out <= 64'b0111111111111111110011000111010101111100010010100111100000000000;    //sigmoid(12.000000) ≈ 0.999994
			8'b11000001: sigmoid_out <= 64'b0111111111111111110011111001010011100101011001111111010000000000;    //sigmoid(12.062500) ≈ 0.999994
			8'b11000010: sigmoid_out <= 64'b0111111111111111110100101000001111011111100110001101110000000000;    //sigmoid(12.125000) ≈ 0.999995
			8'b11000011: sigmoid_out <= 64'b0111111111111111110101010100010101011010000011110110100000000000;    //sigmoid(12.187500) ≈ 0.999995
			8'b11000100: sigmoid_out <= 64'b0111111111111111110101111101110000010110011110110100000000000000;    //sigmoid(12.250000) ≈ 0.999995
			8'b11000101: sigmoid_out <= 64'b0111111111111111110110100100101010101011110010101111000000000000;    //sigmoid(12.312500) ≈ 0.999996
			8'b11000110: sigmoid_out <= 64'b0111111111111111110111001001001110001000110000110100000000000000;    //sigmoid(12.375000) ≈ 0.999996
			8'b11000111: sigmoid_out <= 64'b0111111111111111110111101011100011110110011011011111110000000000;    //sigmoid(12.437500) ≈ 0.999996
			8'b11001000: sigmoid_out <= 64'b0111111111111111111000001011110100011010011000110010010000000000;    //sigmoid(12.500000) ≈ 0.999996
			8'b11001001: sigmoid_out <= 64'b0111111111111111111000101010000111111000111011101010000000000000;    //sigmoid(12.562500) ≈ 0.999996
			8'b11001010: sigmoid_out <= 64'b0111111111111111111001000110100101110111000101001011010000000000;    //sigmoid(12.625000) ≈ 0.999997
			8'b11001011: sigmoid_out <= 64'b0111111111111111111001100001010101011100011101110001100000000000;    //sigmoid(12.687500) ≈ 0.999997
			8'b11001100: sigmoid_out <= 64'b0111111111111111111001111010011101010101000111001100100000000000;    //sigmoid(12.750000) ≈ 0.999997
			8'b11001101: sigmoid_out <= 64'b0111111111111111111010010010000011110011000111100000100000000000;    //sigmoid(12.812500) ≈ 0.999997
			8'b11001110: sigmoid_out <= 64'b0111111111111111111010101000001110110000001101101011010000000000;    //sigmoid(12.875000) ≈ 0.999997
			8'b11001111: sigmoid_out <= 64'b0111111111111111111010111101000011101111010000000000000000000000;    //sigmoid(12.937500) ≈ 0.999998
			8'b11010000: sigmoid_out <= 64'b0111111111111111111011010000100111111101100100110111000000000000;    //sigmoid(13.000000) ≈ 0.999998
			8'b11010001: sigmoid_out <= 64'b0111111111111111111011100011000000010100010110000101110000000000;    //sigmoid(13.062500) ≈ 0.999998
			8'b11010010: sigmoid_out <= 64'b0111111111111111111011110100010001011001101111010000110000000000;    //sigmoid(13.125000) ≈ 0.999998
			8'b11010011: sigmoid_out <= 64'b0111111111111111111100000100011111100010000111010000000000000000;    //sigmoid(13.187500) ≈ 0.999998
			8'b11010100: sigmoid_out <= 64'b0111111111111111111100010011101110110001000101011000100000000000;    //sigmoid(13.250000) ≈ 0.999998
			8'b11010101: sigmoid_out <= 64'b0111111111111111111100100010000010111010100010010010100000000000;    //sigmoid(13.312500) ≈ 0.999998
			8'b11010110: sigmoid_out <= 64'b0111111111111111111100101111011111100011100100111101100000000000;    //sigmoid(13.375000) ≈ 0.999998
			8'b11010111: sigmoid_out <= 64'b0111111111111111111100111100001000000011011100000001010000000000;    //sigmoid(13.437500) ≈ 0.999999
			8'b11011000: sigmoid_out <= 64'b0111111111111111111101000111111111100100010011100000110000000000;    //sigmoid(13.500000) ≈ 0.999999
			8'b11011001: sigmoid_out <= 64'b0111111111111111111101010011001001000100000111100001100000000000;    //sigmoid(13.562500) ≈ 0.999999
			8'b11011010: sigmoid_out <= 64'b0111111111111111111101011101100111010101010011100111010000000000;    //sigmoid(13.625000) ≈ 0.999999
			8'b11011011: sigmoid_out <= 64'b0111111111111111111101100111011100111111011111100000010000000000;    //sigmoid(13.687500) ≈ 0.999999
			8'b11011100: sigmoid_out <= 64'b0111111111111111111101110000101100100000001000111100000000000000;    //sigmoid(13.750000) ≈ 0.999999
			8'b11011101: sigmoid_out <= 64'b0111111111111111111101111001011000001011001011000111000000000000;    //sigmoid(13.812500) ≈ 0.999999
			8'b11011110: sigmoid_out <= 64'b0111111111111111111110000001100010001011100011100111010000000000;    //sigmoid(13.875000) ≈ 0.999999
			8'b11011111: sigmoid_out <= 64'b0111111111111111111110001001001100100011110101001100110000000000;    //sigmoid(13.937500) ≈ 0.999999
			8'b11100000: sigmoid_out <= 64'b0111111111111111111110010000011001001110101000011110000000000000;    //sigmoid(14.000000) ≈ 0.999999
			8'b11100001: sigmoid_out <= 64'b0111111111111111111110010111001001111111001010011110100000000000;    //sigmoid(14.062500) ≈ 0.999999
			8'b11100010: sigmoid_out <= 64'b0111111111111111111110011101100000100001101001100100100000000000;    //sigmoid(14.125000) ≈ 0.999999
			8'b11100011: sigmoid_out <= 64'b0111111111111111111110100011011110011011110000011110000000000000;    //sigmoid(14.187500) ≈ 0.999999
			8'b11100100: sigmoid_out <= 64'b0111111111111111111110101001000101001100111111101001110000000000;    //sigmoid(14.250000) ≈ 0.999999
			8'b11100101: sigmoid_out <= 64'b0111111111111111111110101110010110001111000101010010100000000000;    //sigmoid(14.312500) ≈ 0.999999
			8'b11100110: sigmoid_out <= 64'b0111111111111111111110110011010010110110010011101000000000000000;    //sigmoid(14.375000) ≈ 0.999999
			8'b11100111: sigmoid_out <= 64'b0111111111111111111110110111111100010001110110000110000000000000;    //sigmoid(14.437500) ≈ 0.999999
			8'b11101000: sigmoid_out <= 64'b0111111111111111111110111100010011101100000101001000010000000000;    //sigmoid(14.500000) ≈ 0.999999
			8'b11101001: sigmoid_out <= 64'b0111111111111111111111000000011010001010111000101110000000000000;    //sigmoid(14.562500) ≈ 1.000000
			8'b11101010: sigmoid_out <= 64'b0111111111111111111111000100010000101111111001111011000000000000;    //sigmoid(14.625000) ≈ 1.000000
			8'b11101011: sigmoid_out <= 64'b0111111111111111111111000111111000011000110011010001010000000000;    //sigmoid(14.687500) ≈ 1.000000
			8'b11101100: sigmoid_out <= 64'b0111111111111111111111001011010001111111100000001011100000000000;    //sigmoid(14.750000) ≈ 1.000000
			8'b11101101: sigmoid_out <= 64'b0111111111111111111111001110011110011010011011011101000000000000;    //sigmoid(14.812500) ≈ 1.000000
			8'b11101110: sigmoid_out <= 64'b0111111111111111111111010001011110011100101100111000100000000000;    //sigmoid(14.875000) ≈ 1.000000
			8'b11101111: sigmoid_out <= 64'b0111111111111111111111010100010010110110010110000001010000000000;    //sigmoid(14.937500) ≈ 1.000000
			8'b11110000: sigmoid_out <= 64'b0111111111111111111111010110111100010100011110001110010000000000;    //sigmoid(15.000000) ≈ 1.000000
			8'b11110001: sigmoid_out <= 64'b0111111111111111111111011001011011100001011101111001100000000000;    //sigmoid(15.062500) ≈ 1.000000
			8'b11110010: sigmoid_out <= 64'b0111111111111111111111011011110001000101001001000111000000000000;    //sigmoid(15.125000) ≈ 1.000000
			8'b11110011: sigmoid_out <= 64'b0111111111111111111111011101111101100100111001100011110000000000;    //sigmoid(15.187500) ≈ 1.000000
			8'b11110100: sigmoid_out <= 64'b0111111111111111111111100000000001100011110111111010010000000000;    //sigmoid(15.250000) ≈ 1.000000
			8'b11110101: sigmoid_out <= 64'b0111111111111111111111100001111101100011000100100110010000000000;    //sigmoid(15.312500) ≈ 1.000000
			8'b11110110: sigmoid_out <= 64'b0111111111111111111111100011110010000001100000000100000000000000;    //sigmoid(15.375000) ≈ 1.000000
			8'b11110111: sigmoid_out <= 64'b0111111111111111111111100101011111011100010010100000010000000000;    //sigmoid(15.437500) ≈ 1.000000
			8'b11111000: sigmoid_out <= 64'b0111111111111111111111100111000110001110110011001101000000000000;    //sigmoid(15.500000) ≈ 1.000000
			8'b11111001: sigmoid_out <= 64'b0111111111111111111111101000100110110010101111010100000000000000;    //sigmoid(15.562500) ≈ 1.000000
			8'b11111010: sigmoid_out <= 64'b0111111111111111111111101010000001100000010000010100010000000000;    //sigmoid(15.625000) ≈ 1.000000
			8'b11111011: sigmoid_out <= 64'b0111111111111111111111101011010110101110000010000101010000000000;    //sigmoid(15.687500) ≈ 1.000000
			8'b11111100: sigmoid_out <= 64'b0111111111111111111111101100100110110001011000011110000000000000;    //sigmoid(15.750000) ≈ 1.000000
			8'b11111101: sigmoid_out <= 64'b0111111111111111111111101101110001111110010100110000000000000000;    //sigmoid(15.812500) ≈ 1.000000
			8'b11111110: sigmoid_out <= 64'b0111111111111111111111101110111000100111101010100011000000000000;    //sigmoid(15.875000) ≈ 1.000000
			8'b11111111: sigmoid_out <= 64'b0111111111111111111111101111111010111111000100100011110000000000;    //sigmoid(15.937500) ≈ 1.000000

        endcase
    end
endmodule