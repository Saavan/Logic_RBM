//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
//
// Create Date: 2019-07-01 16:08:17.141783
// Design Name: vanilla
// Module Name: sigmoidLUT_in8b4p_out16b15p
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 8 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
//
// Additional Comments: Generated by LUT_generator_sigmoid.py
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_in8b4p_out16b15p #(
    parameter PRECISION_INPUT_BITS = 8,
    parameter PRECISION_OUTPUT_BITS = 16
)(
    input[PRECISION_INPUT_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_OUTPUT_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			8'b00000000: sigmoid_out <= 16'b0100000000000000;    //sigmoid(0.000000) ≈ 0.500000
			8'b00000001: sigmoid_out <= 16'b0100001000000000;    //sigmoid(0.062500) ≈ 0.515625
			8'b00000010: sigmoid_out <= 16'b0100001111111111;    //sigmoid(0.125000) ≈ 0.531219
			8'b00000011: sigmoid_out <= 16'b0100010111111100;    //sigmoid(0.187500) ≈ 0.546753
			8'b00000100: sigmoid_out <= 16'b0100011111110101;    //sigmoid(0.250000) ≈ 0.562164
			8'b00000101: sigmoid_out <= 16'b0100100111101011;    //sigmoid(0.312500) ≈ 0.577484
			8'b00000110: sigmoid_out <= 16'b0100101111011100;    //sigmoid(0.375000) ≈ 0.592651
			8'b00000111: sigmoid_out <= 16'b0100110111001000;    //sigmoid(0.437500) ≈ 0.607666
			8'b00001000: sigmoid_out <= 16'b0100111110101101;    //sigmoid(0.500000) ≈ 0.622467
			8'b00001001: sigmoid_out <= 16'b0101000110001010;    //sigmoid(0.562500) ≈ 0.637024
			8'b00001010: sigmoid_out <= 16'b0101001101100000;    //sigmoid(0.625000) ≈ 0.651367
			8'b00001011: sigmoid_out <= 16'b0101010100101100;    //sigmoid(0.687500) ≈ 0.665405
			8'b00001100: sigmoid_out <= 16'b0101011011101111;    //sigmoid(0.750000) ≈ 0.679169
			8'b00001101: sigmoid_out <= 16'b0101100010101000;    //sigmoid(0.812500) ≈ 0.692627
			8'b00001110: sigmoid_out <= 16'b0101101001010111;    //sigmoid(0.875000) ≈ 0.705780
			8'b00001111: sigmoid_out <= 16'b0101101111111011;    //sigmoid(0.937500) ≈ 0.718597
			8'b00010000: sigmoid_out <= 16'b0101110110010011;    //sigmoid(1.000000) ≈ 0.731049
			8'b00010001: sigmoid_out <= 16'b0101111100100000;    //sigmoid(1.062500) ≈ 0.743164
			8'b00010010: sigmoid_out <= 16'b0110000010100001;    //sigmoid(1.125000) ≈ 0.754913
			8'b00010011: sigmoid_out <= 16'b0110001000010110;    //sigmoid(1.187500) ≈ 0.766296
			8'b00010100: sigmoid_out <= 16'b0110001101111111;    //sigmoid(1.250000) ≈ 0.777313
			8'b00010101: sigmoid_out <= 16'b0110010011011011;    //sigmoid(1.312500) ≈ 0.787933
			8'b00010110: sigmoid_out <= 16'b0110011000101011;    //sigmoid(1.375000) ≈ 0.798187
			8'b00010111: sigmoid_out <= 16'b0110011101101111;    //sigmoid(1.437500) ≈ 0.808075
			8'b00011000: sigmoid_out <= 16'b0110100010100110;    //sigmoid(1.500000) ≈ 0.817566
			8'b00011001: sigmoid_out <= 16'b0110100111010010;    //sigmoid(1.562500) ≈ 0.826721
			8'b00011010: sigmoid_out <= 16'b0110101011110001;    //sigmoid(1.625000) ≈ 0.835480
			8'b00011011: sigmoid_out <= 16'b0110110000000101;    //sigmoid(1.687500) ≈ 0.843903
			8'b00011100: sigmoid_out <= 16'b0110110100001101;    //sigmoid(1.750000) ≈ 0.851959
			8'b00011101: sigmoid_out <= 16'b0110111000001001;    //sigmoid(1.812500) ≈ 0.859650
			8'b00011110: sigmoid_out <= 16'b0110111011111011;    //sigmoid(1.875000) ≈ 0.867035
			8'b00011111: sigmoid_out <= 16'b0110111111100010;    //sigmoid(1.937500) ≈ 0.874084
			8'b00100000: sigmoid_out <= 16'b0111000010111110;    //sigmoid(2.000000) ≈ 0.880798
			8'b00100001: sigmoid_out <= 16'b0111000110010000;    //sigmoid(2.062500) ≈ 0.887207
			8'b00100010: sigmoid_out <= 16'b0111001001011000;    //sigmoid(2.125000) ≈ 0.893311
			8'b00100011: sigmoid_out <= 16'b0111001100010110;    //sigmoid(2.187500) ≈ 0.899109
			8'b00100100: sigmoid_out <= 16'b0111001111001100;    //sigmoid(2.250000) ≈ 0.904663
			8'b00100101: sigmoid_out <= 16'b0111010001111000;    //sigmoid(2.312500) ≈ 0.909912
			8'b00100110: sigmoid_out <= 16'b0111010100011011;    //sigmoid(2.375000) ≈ 0.914886
			8'b00100111: sigmoid_out <= 16'b0111010110110111;    //sigmoid(2.437500) ≈ 0.919647
			8'b00101000: sigmoid_out <= 16'b0111011001001010;    //sigmoid(2.500000) ≈ 0.924133
			8'b00101001: sigmoid_out <= 16'b0111011011010110;    //sigmoid(2.562500) ≈ 0.928406
			8'b00101010: sigmoid_out <= 16'b0111011101011011;    //sigmoid(2.625000) ≈ 0.932465
			8'b00101011: sigmoid_out <= 16'b0111011111011000;    //sigmoid(2.687500) ≈ 0.936279
			8'b00101100: sigmoid_out <= 16'b0111100001001111;    //sigmoid(2.750000) ≈ 0.939911
			8'b00101101: sigmoid_out <= 16'b0111100011000000;    //sigmoid(2.812500) ≈ 0.943359
			8'b00101110: sigmoid_out <= 16'b0111100100101010;    //sigmoid(2.875000) ≈ 0.946594
			8'b00101111: sigmoid_out <= 16'b0111100110001111;    //sigmoid(2.937500) ≈ 0.949677
			8'b00110000: sigmoid_out <= 16'b0111100111101110;    //sigmoid(3.000000) ≈ 0.952576
			8'b00110001: sigmoid_out <= 16'b0111101001001000;    //sigmoid(3.062500) ≈ 0.955322
			8'b00110010: sigmoid_out <= 16'b0111101010011101;    //sigmoid(3.125000) ≈ 0.957916
			8'b00110011: sigmoid_out <= 16'b0111101011101101;    //sigmoid(3.187500) ≈ 0.960358
			8'b00110100: sigmoid_out <= 16'b0111101100111001;    //sigmoid(3.250000) ≈ 0.962677
			8'b00110101: sigmoid_out <= 16'b0111101110000000;    //sigmoid(3.312500) ≈ 0.964844
			8'b00110110: sigmoid_out <= 16'b0111101111000100;    //sigmoid(3.375000) ≈ 0.966919
			8'b00110111: sigmoid_out <= 16'b0111110000000011;    //sigmoid(3.437500) ≈ 0.968842
			8'b00111000: sigmoid_out <= 16'b0111110000111111;    //sigmoid(3.500000) ≈ 0.970673
			8'b00111001: sigmoid_out <= 16'b0111110001111000;    //sigmoid(3.562500) ≈ 0.972412
			8'b00111010: sigmoid_out <= 16'b0111110010101101;    //sigmoid(3.625000) ≈ 0.974030
			8'b00111011: sigmoid_out <= 16'b0111110011100000;    //sigmoid(3.687500) ≈ 0.975586
			8'b00111100: sigmoid_out <= 16'b0111110100001111;    //sigmoid(3.750000) ≈ 0.977020
			8'b00111101: sigmoid_out <= 16'b0111110100111100;    //sigmoid(3.812500) ≈ 0.978394
			8'b00111110: sigmoid_out <= 16'b0111110101100110;    //sigmoid(3.875000) ≈ 0.979675
			8'b00111111: sigmoid_out <= 16'b0111110110001101;    //sigmoid(3.937500) ≈ 0.980865
			8'b01000000: sigmoid_out <= 16'b0111110110110011;    //sigmoid(4.000000) ≈ 0.982025
			8'b01000001: sigmoid_out <= 16'b0111110111010110;    //sigmoid(4.062500) ≈ 0.983093
			8'b01000010: sigmoid_out <= 16'b0111110111110111;    //sigmoid(4.125000) ≈ 0.984100
			8'b01000011: sigmoid_out <= 16'b0111111000010110;    //sigmoid(4.187500) ≈ 0.985046
			8'b01000100: sigmoid_out <= 16'b0111111000110011;    //sigmoid(4.250000) ≈ 0.985931
			8'b01000101: sigmoid_out <= 16'b0111111001001111;    //sigmoid(4.312500) ≈ 0.986786
			8'b01000110: sigmoid_out <= 16'b0111111001101001;    //sigmoid(4.375000) ≈ 0.987579
			8'b01000111: sigmoid_out <= 16'b0111111010000001;    //sigmoid(4.437500) ≈ 0.988312
			8'b01001000: sigmoid_out <= 16'b0111111010011000;    //sigmoid(4.500000) ≈ 0.989014
			8'b01001001: sigmoid_out <= 16'b0111111010101110;    //sigmoid(4.562500) ≈ 0.989685
			8'b01001010: sigmoid_out <= 16'b0111111011000010;    //sigmoid(4.625000) ≈ 0.990295
			8'b01001011: sigmoid_out <= 16'b0111111011010101;    //sigmoid(4.687500) ≈ 0.990875
			8'b01001100: sigmoid_out <= 16'b0111111011100111;    //sigmoid(4.750000) ≈ 0.991425
			8'b01001101: sigmoid_out <= 16'b0111111011111000;    //sigmoid(4.812500) ≈ 0.991943
			8'b01001110: sigmoid_out <= 16'b0111111100001000;    //sigmoid(4.875000) ≈ 0.992432
			8'b01001111: sigmoid_out <= 16'b0111111100010111;    //sigmoid(4.937500) ≈ 0.992889
			8'b01010000: sigmoid_out <= 16'b0111111100100101;    //sigmoid(5.000000) ≈ 0.993317
			8'b01010001: sigmoid_out <= 16'b0111111100110010;    //sigmoid(5.062500) ≈ 0.993713
			8'b01010010: sigmoid_out <= 16'b0111111100111110;    //sigmoid(5.125000) ≈ 0.994080
			8'b01010011: sigmoid_out <= 16'b0111111101001010;    //sigmoid(5.187500) ≈ 0.994446
			8'b01010100: sigmoid_out <= 16'b0111111101010101;    //sigmoid(5.250000) ≈ 0.994781
			8'b01010101: sigmoid_out <= 16'b0111111101011111;    //sigmoid(5.312500) ≈ 0.995087
			8'b01010110: sigmoid_out <= 16'b0111111101101001;    //sigmoid(5.375000) ≈ 0.995392
			8'b01010111: sigmoid_out <= 16'b0111111101110010;    //sigmoid(5.437500) ≈ 0.995667
			8'b01011000: sigmoid_out <= 16'b0111111101111011;    //sigmoid(5.500000) ≈ 0.995941
			8'b01011001: sigmoid_out <= 16'b0111111110000011;    //sigmoid(5.562500) ≈ 0.996185
			8'b01011010: sigmoid_out <= 16'b0111111110001010;    //sigmoid(5.625000) ≈ 0.996399
			8'b01011011: sigmoid_out <= 16'b0111111110010001;    //sigmoid(5.687500) ≈ 0.996613
			8'b01011100: sigmoid_out <= 16'b0111111110011000;    //sigmoid(5.750000) ≈ 0.996826
			8'b01011101: sigmoid_out <= 16'b0111111110011110;    //sigmoid(5.812500) ≈ 0.997009
			8'b01011110: sigmoid_out <= 16'b0111111110100100;    //sigmoid(5.875000) ≈ 0.997192
			8'b01011111: sigmoid_out <= 16'b0111111110101010;    //sigmoid(5.937500) ≈ 0.997375
			8'b01100000: sigmoid_out <= 16'b0111111110101111;    //sigmoid(6.000000) ≈ 0.997528
			8'b01100001: sigmoid_out <= 16'b0111111110110100;    //sigmoid(6.062500) ≈ 0.997681
			8'b01100010: sigmoid_out <= 16'b0111111110111000;    //sigmoid(6.125000) ≈ 0.997803
			8'b01100011: sigmoid_out <= 16'b0111111110111101;    //sigmoid(6.187500) ≈ 0.997955
			8'b01100100: sigmoid_out <= 16'b0111111111000001;    //sigmoid(6.250000) ≈ 0.998077
			8'b01100101: sigmoid_out <= 16'b0111111111000101;    //sigmoid(6.312500) ≈ 0.998199
			8'b01100110: sigmoid_out <= 16'b0111111111001000;    //sigmoid(6.375000) ≈ 0.998291
			8'b01100111: sigmoid_out <= 16'b0111111111001100;    //sigmoid(6.437500) ≈ 0.998413
			8'b01101000: sigmoid_out <= 16'b0111111111001111;    //sigmoid(6.500000) ≈ 0.998505
			8'b01101001: sigmoid_out <= 16'b0111111111010010;    //sigmoid(6.562500) ≈ 0.998596
			8'b01101010: sigmoid_out <= 16'b0111111111010101;    //sigmoid(6.625000) ≈ 0.998688
			8'b01101011: sigmoid_out <= 16'b0111111111010111;    //sigmoid(6.687500) ≈ 0.998749
			8'b01101100: sigmoid_out <= 16'b0111111111011010;    //sigmoid(6.750000) ≈ 0.998840
			8'b01101101: sigmoid_out <= 16'b0111111111011100;    //sigmoid(6.812500) ≈ 0.998901
			8'b01101110: sigmoid_out <= 16'b0111111111011110;    //sigmoid(6.875000) ≈ 0.998962
			8'b01101111: sigmoid_out <= 16'b0111111111100000;    //sigmoid(6.937500) ≈ 0.999023
			8'b01110000: sigmoid_out <= 16'b0111111111100010;    //sigmoid(7.000000) ≈ 0.999084
			8'b01110001: sigmoid_out <= 16'b0111111111100100;    //sigmoid(7.062500) ≈ 0.999146
			8'b01110010: sigmoid_out <= 16'b0111111111100110;    //sigmoid(7.125000) ≈ 0.999207
			8'b01110011: sigmoid_out <= 16'b0111111111100111;    //sigmoid(7.187500) ≈ 0.999237
			8'b01110100: sigmoid_out <= 16'b0111111111101001;    //sigmoid(7.250000) ≈ 0.999298
			8'b01110101: sigmoid_out <= 16'b0111111111101010;    //sigmoid(7.312500) ≈ 0.999329
			8'b01110110: sigmoid_out <= 16'b0111111111101011;    //sigmoid(7.375000) ≈ 0.999359
			8'b01110111: sigmoid_out <= 16'b0111111111101101;    //sigmoid(7.437500) ≈ 0.999420
			8'b01111000: sigmoid_out <= 16'b0111111111101110;    //sigmoid(7.500000) ≈ 0.999451
			8'b01111001: sigmoid_out <= 16'b0111111111101111;    //sigmoid(7.562500) ≈ 0.999481
			8'b01111010: sigmoid_out <= 16'b0111111111110000;    //sigmoid(7.625000) ≈ 0.999512
			8'b01111011: sigmoid_out <= 16'b0111111111110001;    //sigmoid(7.687500) ≈ 0.999542
			8'b01111100: sigmoid_out <= 16'b0111111111110010;    //sigmoid(7.750000) ≈ 0.999573
			8'b01111101: sigmoid_out <= 16'b0111111111110011;    //sigmoid(7.812500) ≈ 0.999603
			8'b01111110: sigmoid_out <= 16'b0111111111110100;    //sigmoid(7.875000) ≈ 0.999634
			8'b01111111: sigmoid_out <= 16'b0111111111110100;    //sigmoid(7.937500) ≈ 0.999634
			8'b10000000: sigmoid_out <= 16'b0111111111110101;    //sigmoid(8.000000) ≈ 0.999664
			8'b10000001: sigmoid_out <= 16'b0111111111110110;    //sigmoid(8.062500) ≈ 0.999695
			8'b10000010: sigmoid_out <= 16'b0111111111110110;    //sigmoid(8.125000) ≈ 0.999695
			8'b10000011: sigmoid_out <= 16'b0111111111110111;    //sigmoid(8.187500) ≈ 0.999725
			8'b10000100: sigmoid_out <= 16'b0111111111110111;    //sigmoid(8.250000) ≈ 0.999725
			8'b10000101: sigmoid_out <= 16'b0111111111111000;    //sigmoid(8.312500) ≈ 0.999756
			8'b10000110: sigmoid_out <= 16'b0111111111111000;    //sigmoid(8.375000) ≈ 0.999756
			8'b10000111: sigmoid_out <= 16'b0111111111111001;    //sigmoid(8.437500) ≈ 0.999786
			8'b10001000: sigmoid_out <= 16'b0111111111111001;    //sigmoid(8.500000) ≈ 0.999786
			8'b10001001: sigmoid_out <= 16'b0111111111111010;    //sigmoid(8.562500) ≈ 0.999817
			8'b10001010: sigmoid_out <= 16'b0111111111111010;    //sigmoid(8.625000) ≈ 0.999817
			8'b10001011: sigmoid_out <= 16'b0111111111111010;    //sigmoid(8.687500) ≈ 0.999817
			8'b10001100: sigmoid_out <= 16'b0111111111111011;    //sigmoid(8.750000) ≈ 0.999847
			8'b10001101: sigmoid_out <= 16'b0111111111111011;    //sigmoid(8.812500) ≈ 0.999847
			8'b10001110: sigmoid_out <= 16'b0111111111111011;    //sigmoid(8.875000) ≈ 0.999847
			8'b10001111: sigmoid_out <= 16'b0111111111111100;    //sigmoid(8.937500) ≈ 0.999878
			8'b10010000: sigmoid_out <= 16'b0111111111111100;    //sigmoid(9.000000) ≈ 0.999878
			8'b10010001: sigmoid_out <= 16'b0111111111111100;    //sigmoid(9.062500) ≈ 0.999878
			8'b10010010: sigmoid_out <= 16'b0111111111111100;    //sigmoid(9.125000) ≈ 0.999878
			8'b10010011: sigmoid_out <= 16'b0111111111111101;    //sigmoid(9.187500) ≈ 0.999908
			8'b10010100: sigmoid_out <= 16'b0111111111111101;    //sigmoid(9.250000) ≈ 0.999908
			8'b10010101: sigmoid_out <= 16'b0111111111111101;    //sigmoid(9.312500) ≈ 0.999908
			8'b10010110: sigmoid_out <= 16'b0111111111111101;    //sigmoid(9.375000) ≈ 0.999908
			8'b10010111: sigmoid_out <= 16'b0111111111111101;    //sigmoid(9.437500) ≈ 0.999908
			8'b10011000: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.500000) ≈ 0.999939
			8'b10011001: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.562500) ≈ 0.999939
			8'b10011010: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.625000) ≈ 0.999939
			8'b10011011: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.687500) ≈ 0.999939
			8'b10011100: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.750000) ≈ 0.999939
			8'b10011101: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.812500) ≈ 0.999939
			8'b10011110: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.875000) ≈ 0.999939
			8'b10011111: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.937500) ≈ 0.999939
			8'b10100000: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.000000) ≈ 0.999969
			8'b10100001: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.062500) ≈ 0.999969
			8'b10100010: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.125000) ≈ 0.999969
			8'b10100011: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.187500) ≈ 0.999969
			8'b10100100: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.250000) ≈ 0.999969
			8'b10100101: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.312500) ≈ 0.999969
			8'b10100110: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.375000) ≈ 0.999969
			8'b10100111: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.437500) ≈ 0.999969
			8'b10101000: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.500000) ≈ 0.999969
			8'b10101001: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.562500) ≈ 0.999969
			8'b10101010: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.625000) ≈ 0.999969
			8'b10101011: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.687500) ≈ 0.999969
			8'b10101100: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.750000) ≈ 0.999969
			8'b10101101: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.812500) ≈ 0.999969
			8'b10101110: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.875000) ≈ 0.999969
			8'b10101111: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.937500) ≈ 0.999969
			8'b10110000: sigmoid_out <= 16'b0111111111111111;    //sigmoid(11.000000) ≈ 0.999969
			8'b10110001: sigmoid_out <= 16'b0111111111111111;    //sigmoid(11.062500) ≈ 0.999969
			8'b10110010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.125000) ≈ 1.000000
			8'b10110011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.187500) ≈ 1.000000
			8'b10110100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.250000) ≈ 1.000000
			8'b10110101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.312500) ≈ 1.000000
			8'b10110110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.375000) ≈ 1.000000
			8'b10110111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.437500) ≈ 1.000000
			8'b10111000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.500000) ≈ 1.000000
			8'b10111001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.562500) ≈ 1.000000
			8'b10111010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.625000) ≈ 1.000000
			8'b10111011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.687500) ≈ 1.000000
			8'b10111100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.750000) ≈ 1.000000
			8'b10111101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.812500) ≈ 1.000000
			8'b10111110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.875000) ≈ 1.000000
			8'b10111111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.937500) ≈ 1.000000
			8'b11000000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.000000) ≈ 1.000000
			8'b11000001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.062500) ≈ 1.000000
			8'b11000010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.125000) ≈ 1.000000
			8'b11000011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.187500) ≈ 1.000000
			8'b11000100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.250000) ≈ 1.000000
			8'b11000101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.312500) ≈ 1.000000
			8'b11000110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.375000) ≈ 1.000000
			8'b11000111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.437500) ≈ 1.000000
			8'b11001000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.500000) ≈ 1.000000
			8'b11001001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.562500) ≈ 1.000000
			8'b11001010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.625000) ≈ 1.000000
			8'b11001011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.687500) ≈ 1.000000
			8'b11001100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.750000) ≈ 1.000000
			8'b11001101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.812500) ≈ 1.000000
			8'b11001110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.875000) ≈ 1.000000
			8'b11001111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.937500) ≈ 1.000000
			8'b11010000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.000000) ≈ 1.000000
			8'b11010001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.062500) ≈ 1.000000
			8'b11010010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.125000) ≈ 1.000000
			8'b11010011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.187500) ≈ 1.000000
			8'b11010100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.250000) ≈ 1.000000
			8'b11010101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.312500) ≈ 1.000000
			8'b11010110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.375000) ≈ 1.000000
			8'b11010111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.437500) ≈ 1.000000
			8'b11011000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.500000) ≈ 1.000000
			8'b11011001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.562500) ≈ 1.000000
			8'b11011010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.625000) ≈ 1.000000
			8'b11011011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.687500) ≈ 1.000000
			8'b11011100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.750000) ≈ 1.000000
			8'b11011101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.812500) ≈ 1.000000
			8'b11011110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.875000) ≈ 1.000000
			8'b11011111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.937500) ≈ 1.000000
			8'b11100000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.000000) ≈ 1.000000
			8'b11100001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.062500) ≈ 1.000000
			8'b11100010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.125000) ≈ 1.000000
			8'b11100011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.187500) ≈ 1.000000
			8'b11100100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.250000) ≈ 1.000000
			8'b11100101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.312500) ≈ 1.000000
			8'b11100110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.375000) ≈ 1.000000
			8'b11100111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.437500) ≈ 1.000000
			8'b11101000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.500000) ≈ 1.000000
			8'b11101001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.562500) ≈ 1.000000
			8'b11101010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.625000) ≈ 1.000000
			8'b11101011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.687500) ≈ 1.000000
			8'b11101100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.750000) ≈ 1.000000
			8'b11101101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.812500) ≈ 1.000000
			8'b11101110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.875000) ≈ 1.000000
			8'b11101111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.937500) ≈ 1.000000
			8'b11110000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.000000) ≈ 1.000000
			8'b11110001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.062500) ≈ 1.000000
			8'b11110010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.125000) ≈ 1.000000
			8'b11110011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.187500) ≈ 1.000000
			8'b11110100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.250000) ≈ 1.000000
			8'b11110101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.312500) ≈ 1.000000
			8'b11110110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.375000) ≈ 1.000000
			8'b11110111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.437500) ≈ 1.000000
			8'b11111000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.500000) ≈ 1.000000
			8'b11111001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.562500) ≈ 1.000000
			8'b11111010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.625000) ≈ 1.000000
			8'b11111011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.687500) ≈ 1.000000
			8'b11111100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.750000) ≈ 1.000000
			8'b11111101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.812500) ≈ 1.000000
			8'b11111110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.875000) ≈ 1.000000
			8'b11111111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.937500) ≈ 1.000000

        endcase
    end
endmodule